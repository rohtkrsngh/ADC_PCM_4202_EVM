

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
o7NuvGpQAnnRMxApyzRmj3y86EJxftHfP8nHdTtUA9nP7kY8XTo46xhJ03zeLvwpBDGM8isk8hNv
oidBVBIBhJBt0AxrbU4T3gF1QuuboRfWYuAOu15ziAPXKQ5JHFqAUA2MpXl1q/v3YuPY7HZCKt0T
zLb+h43rrIKZtMnOc4YTOjvWlAGmt2ayGvNn+z7UbRueJk3VwddXn8oJEIPdsYZpfZJTZGOfUTCo
2PlMLfeHXnCkb7+5xx7BWjz8G0Y3QDXu1k2eldZb/P+fAJx+guZH4H+46KOaOMo/c34BKvj5T0I8
R8Bj9PyC8e21+z8Ft4wMbrHfQMSBGRX4DR+VG675pwUtQCn9gae60bg/faLF5Up5TMV3zhJPdwRM
aN4JDmR/Pcby8reLfu5FAUgQrzL+buNcVi1LYM25hzRvBT96K1Ftv9SRbUte+LLyKHZklGWVcm5+
GRMFH8q+0b4y9+o2mAeGZepNiwZEFFgUoFiHcgpFTWuRan3F3NORUGmsxSIaS2TWf0goYjz5resm
1F8MVTAUjr8LvY1BfQn4lc8flK/FlhVXOirs+GNN6fLiJZcA4ak+ro+CQ/Wbk16uPg89s/gjoMM6
0dq9F809HninokSvBSGDHOWmKqS9gnkpp/OG4ULvdkU5XRpoJcoUQV6EJLnXkIIhoSPclcA4hFOH
SxhyaVH+UTr/aBwbIHOTYl5Tb//bSqa4VjkthttAsGhyTT8kFBnc30X4E3u5fwGgxQ3Qg4rACfwV
HlHO8nXpZCgBUPIuIA0jodeUAm60fsk/FAeH84zk/PJW/wi+xU5mPuHNX5PFs2vK5wALY5NWZ5Dg
ruvYLcxkkTg6geLjpMgYd1Fyk0JUxn3xpzXMYaG0dMMd4zpM0TcyRSf41Ptgz78tMJAeunQzced6
KqBc/UMVou7qTR7WpnnxF01aFXNeuPHLCsiwOt6z6v5UaSABVdWH6jHfPkX0ShND5CobFNh6CpD4
RLZsP8suJODhSYTiN6GF+1RU0yJwR5rk8hbgroKsKHRJlLkGSqjfFrbCwIGr3mCKMLukVlJRPH5R
O4YfDBLz0oAIQbNnOSMcP+o9xps8EQPgVfgBj8ZTBAIxj8Ioq6xGH3lH9hBLSnYxYeeFzXe3VwTf
G+Y6t9puPgSPJxxkL4gHu+omW5Ae7glXEp10pSUFO8Cc4O+jsG1hlM+AnfdrkhC22Ufibgr/uGow
5W4VWWhyRlj9K0X7TvRdjJ2LF0QrNqoCc3ZAtcaoQsgN98zD4LyuRJKSIzu0eeL/aS3hwz4GIiC/
jYCFHcGM9yWApxJ7dUOkm+RX6mhUjz3AkHtpj/X/0vPjBl+k6WJVOHUiwj+QJgMjpC/bjCIhtsvg
aXukHJHDKRaWK1TfBGx87ADhb9g55YYKuBDCvcYQb0KEO+WkvW1MRU556OZQ2GlrlBb/WBQ5nNC5
cD6CmBPlIBrElenpNqXFtMJBsBUapq/R73vsUsWrcco+ILnShWm3hk0JoZyRa3unartop5G5BT/v
dhxd4rabBzrc8i6Io9iIBx+1oTkfwMvRn5s8VfokaK2hwu+8HfF560FR2hRUIrIqF3+D82B5JWpg
c/2LeUTrvkktbFtcNo2JIx4y9xH0UAbSyvn3pUvovF3BZa3wp7257qQq4uygp8G5q7o3lzTyWcyY
f7HObO/yw3HHaqbXwAVdQOD2bcKczqziSWVMwF7FPp5uif0J8S0mnn/krFcopWMwIz2Z6vKWwWdy
/bCi6cVHvJEjIPcHDwko04Ez+ZUg8ra1WYSlzPoUILcA1Wv9ewvNVGW3FeRESGP9uZFZcj3GT7Gm
c3LvLZLmvFsfQFbypNnbrcqWv4F0u5BdmyW/Weqx7fita1q83pTbGxBfZHT0wJlZNGApIlp5V2Nh
rInbOwT4eidL5Oww36uLjAvy9a2dP0tc+RDmmcKh7fJkNEoWqdD6PcaR1Bk5en+9o18AezJeOA4s
z6JTTZfDHomXaaJNiNC3o1hYZeA3cUcgaXejvLutlGHNyelZHo5PM3/DtDe/HFUaBfshpfWwG/Ca
yjAgl2aODcjlNfHWo6oou6T8bblKSmhHAHqBA0yHzXHcvdl04DU+qsq7/n1npPyxYEIwvdAUO8/O
ppVeOACIs9Fss+EDd1QllS8fVcscdnSRQL/19cibTTwwBOV9CQOVc/BvICQUSqXxsW4V3uxeGNWw
EQ1vwEcBN+wel9AZVriocDdZld9gc0jUDFWHeuby5tD1E1nWh2ihfg3OrHjFUliSSYBUvzZK1PHi
oedL3FvhLnOj8p4WX6/LYTBsLoWYO1ECKS/sGpBij9FjV71jc+m09zKWSl88z5kDBFXalI/UznJM
FDgLgB3kEDUYwV54CzPzuqWjAVwfetJYK4AUm7pMh+1UCEhihbnouw48U8HfrurwIqXggG2dessM
/o4rFX1cAooIDGmuvTUZEtQyRJUoc06CU6pJTeTeGPXgYINPJbVJmS1uRMf2130w8I2454Z+Y4o3
05vFnJy+dC4woKaRuhZe9EB9M2gQG74GpIR3rnm5uN7Ubp2Y+BzlaNMG4NXfNb2h5gy86bIVnbxd
Sys7V/+HbpvH/BNLTn6xzUBwZxKFKA2q/OjSO1JVTiX9VvADYK1L7AW1mxovZePTrLFbd/gjZmeI
BL6D5YHawOzDw5eHJDQjQq9yduUhyfI0cdKHlPR6FzYl5eWGOtNxCcxH2oLn0acIo+KKtr+7omMW
UUluYzx3k6KbgIjduFXg5vveMTB26UfCtg+hoxBfW3h1IbIQOZbCr/Sk2r+dgG+oCYvtU2Q+KWMx
TyLnX1Sby3APKof9KB9l8o3EDKSTcqqvCQO8/+AZ7cqlbjtgB9YTK+gR5+ST2qXu7DKNH32fmoVQ
rUdYpzER8JI/Y3r3Rxal7/dlcCbERmtJ3vNcgWKuIeGS9IdQK2ucUP+LwCTIajVDYZejFtzQDrC5
/5MxViDIAbuTGCzmoeE5y4DWfw22Qbat5gskXi/KcK91hAQd6J5hewGQ5txmreDd5ifoPYW4ZCdI
IKhdou0fTO7gdyZOkjeuOb4fochoywc1c5DpXLElrOTLikBGfv5bnZlT09cnUgTbZJoOFu9b+238
QBD/MBoL6Ky36zyQMVrTb/ItoWDQhqbaailzRwkuITCQ38B5esy5d6jbDWpFVaoWesMAYjyLAvDA
AEs41tGM5f1E5t1rO/ozG2eqp/6oPCep0YCSz3Ms+kNhA1byBZiIHTNh94IfHYnXRlFYp1jCtcAn
B3wMYL87RxSNP4zpsyEdXFzyvrARnpqysqKK5ekME+YcwwFxNu72jBRmP8AFUilqgQumzT49kqYF
9FvmX+urBa/FN9bc9CwWh1Jr6vFrSS07sqPfPyM6puzNSb2GecPYduXowEb43dFpCStaxEYxaAN3
mDUsyayIyk5uf6p2VnVt2vz6dXXIFLL7RJLulApVGtYyTraIRUfFz2m1HWX87D+hTOeVVCAaE0ao
kqRfPva/xG9pDarryGheiRpYzOl7ylmsYBHYufbu6bXpqqN+esp+kZD0lBtErS68+bocMSBTTxq4
dM/nQZRhCuWe4eXGN0VW0yCWHWjpYUL7E/4sNtO1wqMJhe02Gr8ZdxtxToGoDlO6zbSBBGgfb5xQ
fmOrueZJPVavCEcoyIB2yILev9KULV/Jm50UryFFevgWkPmd1pFlsc/iL8/GuTjTDZT9DkW+vvAu
c7LPhORccy/Do4FFcn6yp/p15U1vUS8rMU82yOE3q4ts+83D0G3cYrtj/cNDwRgIiPopkfgmTc+G
8TtZ24Hm0Aq1hjsPiIPp6SepYWZpHwUVELJcFj0llmtqkuLlpZ97nA24pY8Rp7TYorW0OxJW6YfY
ZeQH26IA+STYXvLYlrYnoKGovOJKtiVZEBnFvVaqXL06igPLX4e2u9DNO3KJdsONhDKW8jf3kZdu
t7aw4f2b5+a6ImsOdZYIlv7xmm7SRTrKoOBwAKx4D7GpghfLSaqKqixVKvP17bUHV8pfJYBJDLhz
8QpnOSgVIBUxIGom3hFjMn3bM0Xj2ERufsq+xS7hsKJVHvGLMJwLwdAG//Acwbkwu9/R08abNs3A
21OUvrp5X57YIRhAl/0z59OOwH129xId7DeRBpVJBjGjIhDZwysK8CJqVfW6tdCPfDQEyEW+ZeMi
JQ5Rzo9d3mSwFfRt4zJ6rK0MIWTAaAvDkMmzuEY87iR+WO2CkuMnq1WnpEDKjypJZ2fwiV38aFTl
VcOupGrMI8NtSGLczn9V+2uJK+5UtVyXVhVpuI5JSjGWRZxwZnIjWR6vVPMX6Xns1g1/JLrnXmBV
0cruvULSEu+MIxWRMgvDhe2eFkRIpZw5IJNV8+jFA8hhfpGoW9uebd+IYw56gNek4dvcXH6p/bUe
Dbv+NeG4L2EIrrxwz9C3gE4BlCJMSMYuY+FscPl5D+Dq2eVpLQvrQ7FtHh562u8F3fs+j5W0vrWf
BeZFjqbHwwdAu2DMv7NClqcqYSb9i9jW8m7hcW2vtdlPW6IlpT3+5rs4u9qoh/8ZryAIwZXNNjYL
5b104dV6B0QcMJ51nAIMwQ/Gh1BCJamC0sEdxFuH6qtVDjPN9FyaSNapb8G0rdkM1XueNAYqlk0C
ELDvxAfnJxrLZCxKNBJIVq48sDHOAwWnzYhvirEC+3Y1/0HsEZ21VKiy7wFCVY98Vy5jyIFSPgba
xrGMQC4RH3EDSS6MNnBxy5KmYa2WKfkxoGZrE4MK5EWQTJ3cacgX6ALK27N5pCdO2UTfMc9M62s/
JootyVeyRp2ehkt13GDIeJ9WpmTlxz2FkZQbazIoULJOSWBQ8YbO+AdEJI0oldnMprUvYz/0aLAG
N1hqYgcZrqniMyXBSTekEZyUzrGPc2kpPMnCJ1ghrhI6CtZ5H3mG4yUAbl+klVGY+WSy7HqEd6JO
B9oHygwKbmtLhlcex0R7Z3lhjd3qpSRpGJ/So8ugK6fh7aMXesicmXwTn2PUnhdvmPCsdvB8Wc1N
0FPECi3UgVZJ6AaDUaDs32t+GFbEFqz7NUeu+5GCg3eoc/pJvkxLPqs55ynRfHREaqp1cpSbXZ2E
pwlVhEs4R8DwnQQ9QqxtWeAlzOTiDVFyhPL931yjNenPqdm4bFv31czxMzznmrN1O/5cpTFhLTHl
93ubwxDh49Wa2ZDJG4xL9sTHfPkgBUaF5J4Hqwmvsbysl59JYbxabC38+x1nJv0yX/lvOE+IqHWo
5Sp1hv9dz8q5EcNgpirFIzGXQ9ALITZEzJbbDU+pMibFYaX2wcm7mcLwHim1QTq4EPtDYFVDQqJj
BG8U7ne9B4zyAYbj/+Z3KuqGPmem30CO14WQgFbaP00JHk0zsuYLqnw0fxc/ydWhL9K+4hgDq0Gj
tZ4EG7+szSUqZdyyL3SVS/U58yH5JV2BMN+XWt9mvtzOLR+Vqkv0jvUev6FNc3M27igdewpaMGB/
zPbEZHZI8F69KeAaAyJMaZ5k4W6njbhCgS5smcpZ5AxArOHr9EQLB42EsNHhy4FD7LBxd5lxrQWT
dsPnTQQzGGOfOeX6Fg9x9NjGmAVX9VD1QQS7iMXd1wXSLtB9d0p0uWTH7kcypRxJNR0sv02WTB/b
B7TK2NAIEyLljhUNaIiVSvRrQb2nyjYmWKp4y0AFjNp99UXbR8FOA1FMVFRWBEmHuiiHaW2epfCX
jiMKKJz40dGeOWedOhPp+a6UDmTnUAH/iGVQDzmK7qtdOfBd9sQ4WD2Vi5uooDLm15I5kR7XL+Sd
yteqx59ukvjjyyWIZuQtdpy68L0HOw7F1alsgap3mZV/YWDtabSeTOKGSxO8tY4l+j9WfRMZ0fqA
7tPiGhDvsIRNIGnHDIILUvyN9SSPaExG7AyXx2MLVCexyn+C45RBzRa7igHUIx2l9o4cUGufDfm+
76YLBRFSJa6gNaSNqLJZu7eHy5FcCMmWzeqtzpbmjn6mFRaOX/Gv5mstzSqc1yB0C9ht/2RojhnT
U7uT9yWD5RAH3wg4AP1wte3M+pjc64OBrecKyCwpxCDTpDsqHtsbTjj5qTnpOozypjnTyUZLjEpl
4nuzaaslfWSKYuTHyX0gWqRkith9kNfxVxCDEb0vna2jXWgKjsK+T7XavD5fIZYPZnxO8MxzdCzD
LAPJ+UWNcLlZp4wDE/n7+f5AwoLcWrpJOwQRC5du/2u3vobPoFiGl7TQnWXwq7cdlhXCTm4G9xdi
Xfez321cj5q7ErDmW5SIa4Qod+msEcRThnLK9jEs07I03c+Jym2xuwRyk3pJH2eg2h1ksBkoC0vZ
8ONhnHCIH8qFcTvqxiGfPcYK7Lv1ZhsRKyCzEnQMvonU3riw/vNdvmOGzBwlEk93ZR1YbOXJyoSA
S5VNpFbWp4QqsJle9MZBlPmXOaIdB2bGyrFzNCus2FSSmBZFwryhaHnT7zhG9UswZwvBBlyOP9Xe
6BP+9Y3gvhbsxCx3xLypu35GT9cpptwyzWiRZs0oJx7UMxDUEnJke6BNx4DslWPDMK4NyeZdsbPs
oeAURQhWGs751+9/Tx8z/1STko/MIklXJlp9ldcoQMrp7MDjxcPZlZoAWJGHOg4nebsYOrSM9emv
yjkktM/ipR5z8xYtxIJf99jA8m6C243lSAFdVhQL+ibonIv3TVvCaUXNrPzM00OSTHGL86+fOwKU
WWvIp+0kg8zIg932rF7Vrr36GnifVODJSDyyRh1mkQCs0iqkjhvpV3mgG1GQ+payyZy0KVjmWoc8
txN9dBKD8DJd9uKxd7CDWLrmY9aboTlRAtzU4Q7124JtheyEESDQFXmldgZSJdvc4hGVrHfW5rLp
ucTkdaNKDdrq5TkDEx7LnJqdmtdv1coWz8vJ2EBMUqFf1IMZ5NOuyntjsfd8PrA9wf2mDOG598iR
RJC2tMHGdBLxb6EaGIA8S0IbBcSI3LXPVZjNLFe/l+kNLAhjPqGCyCdosaC+fxOroV1SbwjGM/gF
v03y/8B/WCQePRS4qQTQ0XW4Xi/OWNWBS9WYcqquMF/ry1sMjf5jUkB6ANYM47GSk3nntGUJ13Uk
oyC+ujblWk1Z65NWo0ycIASIRKiRpvASyrpiWJkU0w/SrQy60xnbXNodLZz64jwf6ejK3b7FPFUo
0Rf9p6w8UM4aJs6mjm5SZL1PgvvpEhL1cNGV1LfYbrwg+Ng4beWMMPo1viRsRFurqrURlV6c11IR
1+cT1qdnYbd8GHam6moCIkPi26GLSRevKzb6fzyLLyTbEsE1efMSYe0cOaIAuzGxbQj/VY/9ZnJT
0RJ3CRGE23KFkjhDDYgJyXas1mKduR5D3FkxrYWQ0hug7jUEX8tc/+lSCz9aShxEVITRqP2mnsbV
aQ373wPDapEtE8k/BkCGrU2rKJ/8r3V3R3oiJ/OFbGekMIl4d5ltc0LI7nicBr8LEFFcaO5nIrP1
ZVg4YQf+B+t13qcN/1AE86XYiwQwenOrh6EUEEYi7Fi6iy7MmElh3H/F6xA2zPa1Nlts0Ura/7eA
ZhDYIANbJAI7eoLBX+iszRZAYYFl9cd0AdVw5/1vnMsg2q9qpPRWqOFd852AEZQhg3qVqIAd0QEO
OINzCiiR1ZO0bsfCfJcbrWb3KryqJDl/U8L05FY3W8lhNydqusRiW2r3fFN6mvlzX4iIXdQKtPVZ
DJMAmZWdYsr9TM1ne2U7mWBjWlEtsqgJgPm4Y85JPWJwFT1jEa6XEo6CMp33Qt0oKhVXjXCgc0dA
9u5oHxJLJB3HLxkx4fyPnClkzCtW8f0TsMSA0+QTiQ0cI6RxuSle7tf+FZxr+JGXVRbCI8HnEwXZ
ETOF86nb+Ul6rrNKKTV9lniKJqPt4SORRmkr37/l7Ogw4OoyoAbhi7viwgFN9u1S36R9jcL/Ynwa
ouqkZ70r+9dBjclP8G2NB4HgphgtsFvBk23eTElbajeDUxJ6VEUFdxpd6cMO4pZ3pqsKOnWC67Dr
Y8gsx28JBApeUVnwuHLqRFSfZ2CrVcoGRTCxeKv7IGH560CfcTI8erbymoa02BaXeB5/kRIaAOEK
MUf3pz0RLT6pb9ALL5k+7aT8ZqHi2U+eWeKLUjFhkT5sjUXGfPFkWVIpeZwEma6zmyaFqnx2d1l9
KDavWnV98p0e83tG1vOIKo3QYzbpBC6+gHeHFsywOtSLKZ+zZnATrv1nt2y7iNWrxp+x4mlkjUZe
hoMUfR2O2zO7ihr6YQEH9ObwNsjZBzAwWzEXGeXXE2b3rptJpaYckLaQDtJQEccL/daPrlKRwGUH
xCzGj7hpTBzdXl/QXdn2OAYJXhA3iJY9QEtPQIvPOml2osBm5K04F+u1elYyIPiWGXyI66WacIir
La6OVHbwH5VH8lu592f1QO6vZxeRyf377VMfiI9GPlSSKipfipYK4Hon1RxX8/jYT8M2aAeEunbc
ATUUsiRVDa9NohV7ea6SYoWnUEFYnuzkVrfPZxnGe7mMteJtT0c0N6HVadO72iGDvbDrmu7fjptP
xqab5+Oh0tnzPSds8ftT0XvEvTWP2rAJ64Z3IGxyBGIw8y2PhmMdfBLBw4saFuEM4NRl/PLAQKiV
41j+vlktUczyYntkJtBPT1LOpiZy4vo77VObVsPTy3GdgxemEjXdbXRYYXS88yKny/SIHT9fxYfY
jKKjTA4knXPTws61C8XigRpXrPFyyHQojnU2WuehSS8bCi2vvm/7SZ6T0vjO+Q9TJ34CE/T8urlW
98kbMqjnN3LegiJmZTw+GXPLDXPPYTKP+8eqbEk4V12ejtWBWWQCW/jxTaJa4Q7RjYR6VDHQWR/H
OwXLTBIRpZPzYrnQu1ZOepY3YQSl096XCFrNsgtgSQHG0mQBgsGTgqUjBZiwtzH/yIHlAfXpXzgj
HQUz5d0bfZob7Zml/thlIYBd2EWjzm4gE6RcYZ4bm/w9lqfZCFEziuItZ8h+AATdcy8ZbR7XFAND
d2/KUlqfc6I2VgF4boM5nmDUrNw3QrzdUevb/FrSJifZ5mkbrlCvVG5eW4RpCLmcago0d1Lt+nAx
6K6IB8KeE2lzQEwg9KtCPvIwfs1o7p/jkbkS502MdojIU93mkuFi60Rk0xMWFdyZzd1Y5Iny6Z9M
mTq9+YOrAmP2K3Uyx3+w1V9TNSElhwesxOFmIqtUaUA5TTHq7k58sbh3/yLIOyESg7NK4D+lxts0
pvMiNP0CmREfxpPVUa5iwmTxmEVC0d1zUoZiesdga0r2tGL+fmjQ9o0SZJsRyLacu1BmfAkGjvks
nIViHKMM7NEqtiuyjlm4Wg2nVLC8z293oTJ9IiMK/uR5bBFmo3jEpBQZSxyFW4/nks6BFw37PXaA
xlZxJ4MxGcjUzfKJ8u/THBD+pGmrdVhLE+VA9/iT5lConDuRwX+E2+PaqFNHTuP4IfCk6Sd6pSE0
nSIwzVh6PRazk7LR029c5nINJXAPEO489uw364tIeELG6iw89u40Kg0TPPA9NB8go3L3Tg+QHF+C
3lj2DjUq/vIBQXiU98fJjfQ2ZTE6aaByN29rMQ4qJVQasvYXLlAl1dOBcjkllPynBjsWXgVlk486
MPsRo2ctCnWRcto2FpMl6BttmXcUybTnfiwZ6sCLMITsja9bWov37xBrpG1h/x7Moc6tM/L3K2lA
Zhn6ovNpP8iT/dCKO3n5+qbjfTb1Faqk8lFYmhAh6+7e4bQfdUuhX5+73OfyeCTy18Iq5HfkpxGG
5MGpfiliwU/AXGblteaiVTIeNZCkaOXNlygemiZfeRjvw9n1PZEP6ePUq3+r+H7vxb+94NcA4KPd
f55c+ct6YsbHgil0lFrbDG3+gtHge0XFCuZ9PoTLm0nKFuUqLr7M21SYHhfQ8f8+4eA6r8yBSgsx
t1Pf/jDdPJbvn9DIPxsrXKFtCa/YTM0WXIfqiFLFIa/0+uxwIL54ZsGHhGGsCKDpiHbx1fQYiVsG
q16Ce/xhgwTdITXzOFIfIe2MK+0K/9r7RkXSMIF9W4N0Tt7yO9wV9os7LPYSckOlsvPbwFyk0XqM
RB0IUPQgpZpKgn8+pZwOqbYGKp7CADhqS4enN/gRPMJYcDN06y0GHjy/65zrDKuGp/8zt9HSYmCZ
iogsAYNas4KS96qJQu6j6oItWEUjF+XBFTXLLN5cnhWbt79RqQGAmdTnn06Xw4GvjYMliotkt2HT
KSnOQ8H3+ZU6dDWZUSOrg03CRvLG2IidL0oBhh4lwDgIna+ZgpaVT4f02mhJGx37ckl1zp8wh32b
PvfPAEYEqMbwD0knXAT//wGVYCO8sEUakGgEDtijYLeyQW/pZtSYPKl2GFMuEjLLAyjNVMy3wKNZ
hmKWcTvIPeqRRjLNGSg0mX3ZoJ6IE4BYDeDc9fRaGozuMKkA9FfElIsJ66SRndFdVaC71m+Xf0On
kuxq3zgyD9SjHirB+ZdMzqDIXdXt3ziDhNJRIdlAWb5xCwqSr9zt1sa6olR9o6fysK4omlsD+VNB
8yhsnXNRsoH/aVgaYi5SovIWyMCc5k1y7bRRoLmG5p8oTw2VVKf1pnQMel1fuwVvSN9w8dEZPzkm
5h7RyOO8qcNQPo08QB0YSfvjWbhZLlHp1mFFyRDZOOjuND9XhzxTZmL4TC6w+YJzo5/3OOW8uSol
lhi77/Uda8h8MzGG2z8QK6/vAOAzqtshB+2HgKJF7dqo3h2o4JM3E/HQVBc2vrZiYEE2pI4TbFUG
w4oYGjdDZ2MxHCKoGvJ9xJwpes/CP8N7lXQQnMv+lIHgPv2dkSR+2QotMk2HyG0XBQMb+Xo8ns0Q
cOuve/qjmoBfmPZDMjgf6PjqN6IJd4IwPl5naW5r5n5KlwwdfCa0B2EXMJ+xPjjlN5rVd14DXCQM
2AAVzhnn9/1fkaJD2g9lGpUFx5iQ5gJBmt+cCzVwcyHbKKOuVGK9NuErtLhPcsqrXG5FkBh58XsR
tpb94pjFfw5kitYj+kECX+IQzMTmkCr+BnBLaiUVzXUbepr9QtB9oPnfM4EtqM2nN8wWHxd0tqyC
fXPfxFx6wq42UtuliFGJ5X886gJmzMszFZxpN9mi2BJGmTRH/abbyiYzEvJnRkpnsizr2ng2jWg0
lqkjdr8X4sm1JzLrHBtLuqLh2P04i+5kWJ53LOaw6UVbpXocIvhyLu09U0sbwiTIrd5mcQOPZ9ay
ZT0Vw7v/vlcZxfmTJW393ag1mYlOjfVXGdR2nbPR6I38gZLOro1QbDgLircoznBsXux0/xjgjm1o
kcT15jeG0ICE6/M1JPbvlvgianwP+B+g7RwRUo3DgEUQWgWYVkwrQc5CpcbwD6BbWLMlnBKdyq20
pkOF1EZ424K/jKkz6+xSZML7gejczWF+4R7h9O9W24YMLzmN0e5W+Cb8EjKaFQEKDQ7cKPDav5Wv
9kleXECyQkpGch9fiZU0KqA7SVZ+BZ/hGn+2IvA81K5j2kFa2SD69RHncHCS6gWstvDRVmFHaY/u
+KdesDftmYYrYIyYBTz1JRjhIRwQVyjIpLBqpmfmFWkfB0EdpacyhY787VIUS5Xf2ZEFtuqmhhpV
t+v1HRZ6iYKuCo4vbplWBztg/1vTM29ceX5NbqQwLNztyFfzyE3dEjsgDEw3QAzD6EBW/1CuxHQ5
3+A9xR4c5wp4AvkFrc+Ee9iCNsyqOaH0tBaGqWFG4FbW1Ox9nB3+KH/27K4+2s31zdB3jV3GqNi6
VZoQglzzGcjkFrbFRPhNyWLYbSircyJoX6Xfummp1+n3Uvji+sRvLoMXZV+eagZrIRo7JjUOKvFq
s0HyMjW0zn2pD+dugajLN5nuMQtqchxu/Uk28zYo9Gv/OP2xViyYnNi9Cx59zTHLpVr+H7t33Iow
fgG7CDRzxBw5U/ZGgk6UnTzmD3no2GNpK27rw7LT+qGY94pOmAHXl06MoYF9iep7tRDhhEe9VI65
NjAUwwErSjPpmfasgnAlPFBCEIuhZrYfCS+hupgykAFRtq/E3U/jEkFeogSm45gQry6LoRs5dpcE
MRESgDRibFgt/MYVmQ1mtysvUQznxZ6I4G14J21U/9zXZ1uziFwLjHb1HERCwTrMxU7TIPyDyHiO
vfE2jn/j+cBU4kSfCFV/cujO+lOHF7QtbrUal/E2710ccqsknXiodS1QsdJAw7WWC3Ho+V0j2Pef
Wg0CkltIvidAcNQdHH12ttiI8GbPJJTpnZsmHnFbtUqSojJ2O2WSc58FdGzgF8jBRzqsF3stGYSz
LVCRg0/1K6z8ZrJIrJHjIC+k45Shcc32UiBmrfyy4iyR4t+CJD13Rois9IIrymu9i6wEvBnUnXiB
rTzTLLPuJMDL42RgVrXe3bAXBmzyhhIcrnVFbpUlRGFlr8ydUpaJlCmK/sjR+ZaiWn4z2pD+GFPs
cw0xVhUw2YJNUt0177CxrSgYbqFTx8IG+BLCsFSxjr5vztBkTG+kWuJruyYo7R0Us6OaN/BTQS3C
cFSvySLoVjmy1QXvQBKJa7cA0gAr8IzMmIkvTIH/18PwMmI0B6X8eRzxSpLBH7PjV3mYArPPu2wq
0GvJTg7rrZHJaTsEWPSJpzyEK6mVGt+KOT15tB2LrMoGVgd919XdnZVFhQAHTvDKjL6iZkbXCPxc
m6fZcDUp3piNB9CAqrs2bAYCf1n8AmNhfL2lbZbG7raqWGJRmTMDd7gQLVmvhhX8tdJowROJESKO
MkFiwi6/RjT3AfbrEgED47KloTZE8r2ym+VEVIUbVXij82Xg/XUN/Ci2hHlu2pJI1ebagpg8PveF
r0eviAv0btOkPTrOvBUymPfK3MoWmCRueCXx9TZ74aIMD7tf/iXmUFjeX4Oc/J0K7NwFh/XvxEyq
mgRxkfLvV7qLrqTcS7DSiQ0SRDucd1SDWuwfhMJp25+RHeDR904Yq5i5LCw+vz13V4MAcuIZL5NB
64mkcSOpktNpRdX7oOcEujWrSp3x0TYCEq3t3fn3NaI8MEPxuT5w2YkY6bBaK+kh7pgAV0NOgOgo
bM8il6BIe8ReALzwXoR78eF63W5EI5+mzowntaizFPcn8ngmkWcJcQc0r0yWzTO9rlkXdjELRmnG
4XwraiLnoxXOXQXf1iIVp0onRB/3LDp+wAp5dpxFkM9cfP9DeZLEK6tofZNOao3SaQEe3wlFfFQm
RCOjQRWsRraN/1bisBnhblRAPZM6AiR4DGJylMpcj8UIEkeA+gOPnqDB2p02u7Zs4gzHV2p2Aec3
jfZj9rZlUZExfNDIKhsG0p3WdvkPlp0S6B8y7h8YqtD/+js8sM7xqkyIfrfC47eoETleDvPulufN
o80/1B0LIcA6IywUqpYuYcOZV+/yeqQtRBRTE0DSAgS79zLm/N/QKYH/Y+xNxyepzfF4pG7mAsXC
BuH4toh4mbK9RWU/GA21blfm4yLO0M6D3yoY+ByPBLBAkU2h2rQ2llciTp6yQnXUPOhS93+OLwp8
magM4BQ0oXOlXLdWqXwJE/08u8duGF1yR+kOVcmA3nQvJ2gdMQPvuhI7ID2gbob1qoVUnAQCkWmX
wINnI9fSbwDEsrESyLE+vtap41vHqXgfuuXL7bBi5aMTVwiU8+iDDGXli5Tqv2+erdP/VKBxJJwJ
uJp0AoEqKcC/qyRCY13G2J4aAgvJIXD1y+BqQXtCNILZOIsxroPV7xa2YBn6nKlJxQO5HSZ/4rJY
jWZ9wlAXAHf9YfGg0zDGFxgZPU538j+B4U14qhVxvMiG1fg/GheQv3befH3I5SQ2gFWFhJDJYR2B
DblcWdjme+d14I9WNMoBbkIbMKNH4gQoO7lVdhu0EjEuZUbAAy8YJpTHTxS77uYj6WXBJNkhPwQv
tCGqE8+NaxqCU098WyjGxiSsNicLfF2J+pJeYJ3qCaOySg8LPi8BJCw/UNF2kGO6wkxb9ToQ60JE
F/kSoedZr2rnUlXUWKmgIZnIucHwA5PcX2M3UcdYq3VMB/RRzEYCdgYS3hK8QltFdAoYHtZ+DwG3
8bn/IVQnY/IlnGoThSL+O5XNIBvq77PEqKzdf6P2/klKdXaZPTOJ6hhkFQksXl4BewUphA6SnCj1
rq2xVFXc1ObZDqL8tdx7jgtFBV85GQqENRPpDPsMFYMDQpipHWxgdQ9TXHCE1qVGx2GmKLTvf9jf
X73OGadqj0dl0X/v0eNh+QWEQuZk79ski3zm34kB5RM7sOKI2yohuRP0VRbn6ruuSbM6xLnq3JGi
xUeUziAQkPR7367uG17SSuasSxxTBw/e9zu8ZSyBMNdhR4KGX3diKFB9tPekb3d0eSA2tK4S9uOa
Ve74+VnKITpcxKu8AYJDeYl4e567ALIxDDYAxuxLJwRByciZUzwddMqSarufhOAGPSBjFoxe3dqN
NND04+0weZfVY/ZvrsCot8em8rtuGBHNe97KMPGvVycVxRNkPiWeZc0oK/Auj1GcomjkHFiFYa6g
+Z33QwymOMOUr7ZrX6oPHWFC8bFanKq6H3yk/bM/clMCNay3At0GhA/hqgexbMwtBlXCTt8Huwui
hhF0ZsIYKKV0VDfSETCANPW1DYZ57iR8nkbCe62NxRU0APZRx0vu8PbT2NulgQ8azgg0jW6U8TzE
ykJbU7f34r7j+6YNdkC8Ek7pgzGBLWBkCFteb1o4hyRdxXHrDLLVszPs8UI1+xIv16+otfTD/M5B
eBzrRRy5nN/9YLANnukKdJPFCp67WG47/V/obvIEAoC8/p9W7KRLeZxaeQprw5CHKUV120OzNQwk
a4mxB8OWStWuvJJctbayf3oJZOJ+OqElIhSrjHFQWxInDaJZ8gyYCXp+DruebnSvZHcKiWklnsEV
qbJRzMw0fzm8mirpJTs4pEMkxUEUFKf7r0eGQjiUqw8vRjtAhpWobSQzdih9JaXb4NVUFb4UgAGr
bq4jGw6WiYwp+TS+5hmr3Qs5KIjbKmr4Ja/cObyEbF6os/NIRx0ATysjelJzIhgdxnZRQ0Tf88au
yLrLYX1gYqzciBVxw3Vl2BE1Q/CMdo+Ho2M3JA0/yyn6I8pypIUlX00hwNbWDdqYDdotRo+PFh83
LVVkiQ3fYl7rQD/+0r0AtGf/qiyU8AlDh35XBShki1+50gGFHbO74uWFQVFUBU6F+vs7QcRWgNWY
076JBdxO92988kAd4tIr2e6hUxkx0YydbiqVBmNLw9IWQyrwQJNcL7VrqbDD9JQJpXFpPaSE2BSM
EX8rN6xJQY1/8FwHo8Py57YI9tqE74FR93b/ADEZP0FmPTEnX5riPtugmUz9ANRXSMU/UdnhANRs
UK/exa7IY6UkBmZjBq/oyw7Ajzcm7BLQHumhKhbz8Mk0WaKDbRUg09ppXRFcADvST9bxADyzuzTi
fqyx0FLkMc0NsutcQcYjKB9byNaovzrlTbIAE6tKJyYsgdSVy+uLdQDfw+FMzVI204hnH6NckyNm
JDi88u/CUjNdbjVgMu3+cDKezbEV0gssipDfpW4jZdlvx9SrA6UOi41U25nID0uCQFf1vcXt27gw
/gA5lid+7+UBOz4rUl5uOotNSHnNV7NvJ+7X3eHU0cIcJStbaTlQjijwdu1eo5j7K/WINXxzf4Bg
bjuTs10sSBcl8RRHtLUS5dj9mcFqIwQ/QMVW+KW/jbEtOkMZ3z5s1RUY1fg0PBdU/7PR390Vi2e8
99hgvqMz9Cq5o5wz7IX7w5Nol64xvI98T4rQERrK9EBD+lzST61O9eFQfaq6IDX4/oEFCNVtwt+o
JAzwnCedmql/ckHonuVlGCr5NRYGz0JsVSBeGBeYQG+/XeDjaId+MEodS9ULOjq2oe9KSLwBxHlb
Jb/apuzm6zdaeUS8J9nPr2odX1Tg1jqOSA7BhpKHrDy2+4XXpqvbt6vnDWEVpPQwksElSdDGZPsC
ClYJG4rnzHW+qfat0CkgSKxO3xyNZT7QrFvAjFiqLaveyl4JtT+l+k5ySaYdRBvSf74/6HQN7X4r
TRKzwov4n6tN23aRjFs8HQYGIClP+FNEXDZHiotpZLzd9sZHYo1nOogqHJty/NmDhu4Tet/wbtNL
uKMCts2ki+4dECJbtR8ZOVd1WaXFSIY204vaIk8wlBKp4922UHCP1ttb/665/e3EU5u+SG+cz4NM
0Id2WPaOFZh101ykVWxqGiNC7plGewaRj0KA+JnBO3/TWRGBgAqq6wdfZDyLwCKu7VuxI2rfGqSw
kpqtQbjR71K/fyzcB9/PCR4g78++S3gCqG3C0oqHMvrF0RBWORQistccOuzEwvJAMr3x1Yza69t+
rkApbJBkiVFPEWgNY/dT+SMAyW9w+obf6NyePeL2Ngj9eiml/XoM95OIK46rtFI8em1+JvK4ZlJT
vY0Nk8wRfnVvETbwyD+Ks/KwRm/zCjtg99fTHFb2kM/YE3nZw50x8b1cPXr9xbOrviysOmpz7q7r
V5hA7lmvsnecZ1Jd/t3xLLFkaD6GRam0glcbFSGlOY8oHO2IPzTyIIGB1qKKHlmdw60tngWBo6y4
3liPZ6CnQx0VPzKr/TEOD+arKv9XAy3BGSCv//G/9l6ZE0xSx9rmuzTEFw0p3f73+kLzDhSbfC/1
4ZKlNOrr24+hF/4PRvB46RtfOxH+PETmStvcj9XfutWMgRyfNUxv5uGzb+eoxNRdBchIkJ/8MWLG
K3JOzRs3vijXFBImfCLZw0P2Jbe3YBfoEjwhIH8O3DGTZNpPDvaKuPaAOlYP/rCPkuwcnPcGiwRo
61/zqtD6h3vd7ICcJPhwCd7szOYA++3VG22TDpz8DOZE1DWWjoVrxV/67QdwlCls//HtcR4rBToh
74nNT1052tkwkhskXmbABXiQMTKdt3DctYJzuUUgMINP+pZuWn8HX8W+KbKtdsHubVo/xduBX346
HisOWAiJ5MIcUNjO1QYz7tiDMDWc6OSOHGHyiEtqPQ84u06O/BE+E1G9ugcEpcOCT69BiO67HeEL
DFuLChm/yuCVAK08+Pxu+Jm/oYQ5s0RxthUAJ2z5PCiFJoJI3F45Sff5K8hIBCxXr74O9gyr2i9i
mGqdjqR4V8LBHxlzH7c1AGjR0+MIJUUzilWxS9GryY+vh4AGuFpf0p+AMH/AftJdkbRwVJxE52cy
XauQ9m0ikCUMO8PiDEfyTD/P4jehToLFjFRnZT+vQLhFTls0zsQ2d+KilqHPcXwjneYdRtqJYkar
v/tMM5ZE3id6byXiOq2Vh2iXdtQtngSbPZOyBOdZmtTJ8k2CpM/n7jjlErg5e7KdonJy5iF6ght3
97L1Y8vbTsHAC4NtEiVmLy92b9Xe7NnwgpfxM/FAIjkTzjX57rg24gsDVwNjLuudNlm+ptrMDz9i
qWME2MDjQzNPLf8QTqXa/80jm0tv0kBRurtWiz88Ze3CEAk4yxPVn7RKfxonR1d89kFZX/2EKI7p
TAIz0yVjHMfcLjTsLLMNCzMJ0aUkdX4bEdkB2jkH1EFibpH8YMlZ4q3j5vEmtBeZby+XN4zHo2d/
VqgI51g+jy4l/CTXc51eaZyOIXFOXZMRcYXI/x0V7jRGKUb+vtmXlXq6aYYVQBBeGN3xfOMbtGPn
SBJbIiL20uET3v/gTDOEjTKEX/rlskci9Zd8Fm9X3myRHWpDTej+Yedykzj7/OSPWAsAmeBbdOAX
RK9iFDez461uE838IA+ttyssnNHjHhmXiTdBGtVkxCyQb7U82OXFHz0GLJofY3cc9sW8ucuEYyga
+AFK7/NuRkoq7f98//sgs86BsRy80KxgdB38cXzEFoNnQTBsG2LCtn2nXo6/Dfnk/HgcKYG9gS7O
YPed/5/bwqwueyapzynxzMx5HOHlwgD5j2H/SBA1LcPPQJDNbWW84Mps7sVzei4xVLlpBTEpT4Ev
cFsFo2snckoI8Y6AUCW15u3QfbwXE7q0oP19CvGkqdyPR2XWvVa5e/YcuQG1+ibpVpi0GJPN51Yf
2XMBWcTiHRPqLSlT/90kbRVCBFdSU7UtCphDdzRFE2UJ7i5OQ90IJaSkN1MYPA3VSkdl/fKz2ITn
2493XFLEEU4eOG7TU96mtpFZ+ZTarb2LWoO1azAQo4XUDb6eEi5BhPkwD1VgYeCg5xJf+TOhBwub
dxam2I9YPv+KnveMZVg+jjjDYHhLsCN4FRaJ8xG2wg0Md+HE8HUYPfYKYHT4C+1hbHxGIYs1ojcR
eVTSU5ZYc/Xda74XAoWH95YplPE9NniInx2vvD21LwhC/I639h2skulOLdSM/JtQnjt0GoIy32oj
Ro5yEJ7Ni6xg/OPwnnHyALeMUetQ8wp8gbd1g4xtGwBoAhVOIRzGtgAxATRL8dzehwLdmPDFJYQ4
abgHbtwpb976OsrNQUqJademHWZ5qPSFwJm01ZsnobLxETHnEugvHwdmNg1OQNS7TBA26Wn5fxCq
6v4Nhi/N88r9BKpAwVS0BiGL6df7i4XPCN3Z5bQuvXTVDRFcDJutyY5eg7E27d/7BLfPdgkrt3bi
cg9l3OoP1nNGHzNwXYl0dDv4kZgmc6TOILVf9f9RpG8Levuiich26b07rPuSTKDFIgrvpEHy0O76
dia/tTohw6S8qB5+O8xMuEowVyhzaz+34CG0lSH+F60HwjPYFzbyA44WCxspbVfqj3ytTvd+DNgr
T5NUgsjJvrjrEPCWtSM+s12s1BhLSk07mS2/h1phyweS2wNuPwEYtfEgXjhModVkDQ+9fhSjplPL
aw5j5Tg6UR51BFQ4oFkrTgOKx+9Tti2DT6+6H7LJ0pmo2Y5Mky391cRbspa1F8vYY0FkOMhu0taO
GWYGnn0QtXLZIz98DIe4ApR49z92fz5+SdVFc61a+TreV3/LeOp1WvdwoT4j+bi76td7JveBafXu
IDBX9I64W3RajOfG6LPSsSmlzlPB93gDjC3IapHYUsIRAEyYbVpwtwaEorhyLWRLpseNt0FAlTQR
rLmeNvkWqYlwn6il8bh5RuOh3cFkJMMyqVPKJV/zDHgiCUfrOPVAA3oiHSjhoef0iAyh2OWTkNgy
+19jeKwv3jBw8IBK7LESJaPMGeCdfegn6Q++1J1EfiNjl+nBUm6lXHJlVSDxodNg6VrRgdjExluP
2gMpF8JF09brFGWF/o7zSe2MZSx8Sqly879LhxcHD/6aIDYp9RGUdtnvWtvna+hSwdDveury4UHT
m2dUSLefW6XJnARJc2dKXezeMNNP0X25n0aXU3z4a61SH19EN/Bihfi3sST569udERZPRbUFo/b9
jMYZxt3o6B6dgcBgX80JV59KUBRZLQqL13682+O7rJKrWkkG2DU2yO0qr0mB1KGI/cNfVLgpoJNk
Y6Y15WCelVLtx0SVc7J6Y8IRqF9SNd1sE30FH+uQ17xk5F89iVNXMS4RDMQJZRzbRiKaEmmZYQEo
Ai+5x5N3V9MHNx6zQz/3tZVegj9W/+TS/niyRpz6fDx/zssisOz6snTr216nBr/OLphQ8uG+WIEm
R5fGWHKTicyHF4DdtWryHRRoR6bl9h5EtRWQyM01jZt/WmEfQMCeuFMJu9FI12Y+IbUr4AGX6T1N
gPd1oS3so7mc5g5n5+ZvJDJ5S/+c8Ul9/ZXEWk+2hNANkXLdUSTqycgXaF+mWXJXDVEwn5w2eAv3
tIxtCB6TusQjPVI2gLQl3wDlKQCaFHyE9VzuZwYRZj7Uu/SjJcYNdCis7fggkyHpj33hE8Ujp7a6
SDYazThdiCOwz5B0+s+J36uqT2v1aIQcQ4WDKpGJZOVqWk+27LCX5+7AWByfa7cFA1PqiAFWQjnE
diDpFwqEgv0fFHE+VhEDKU657ekUUqj9l0lhyjr5ABFvmldTnkR7HIMhy8McbLZG+CiV3U+BKJKZ
bLJaZzx3M44LuPvWcZykRk2q1z3GTdiCk4BoTVYlyjahAiQq4OxiKYCKOMAJMPQetluhXSTJF8eC
zCsPZJDKRbPOwd01arpFzojEEucwFRoWlaaH+j0o46YHDa6ZWbePzr8zVYhzDks/4WOi85tz/wFu
pMHd4DiOH3ztgKBQvSg2lX6vwptpEoJc3pJ0TeagAfePztCCDPboH5C61YI3Qh4AQ5JU6/JsjkoR
LNHEcTA5Tw5mk1R9ogDPhSjF5qFbQefpTfodMmSCYbq8abmotgt24CmaTBOYEut1oVGy5szdac2X
PwkSvlYw/jEVTkydMGa5jRcuO7eAFk2ueCbs4jmU+vz5ho6dGgWftmf7OYENtRtyctHd25yeC0pp
Lxr6pPuyOEDw2xxLHYVglI/OawjguQMgBnSoyM0nlQ9GnVLqZCeLTGB1oQyjy1a4UxjX3FUQ+8kT
+pVWxRsYDEsVdt5aJaOnuOlYxnwNiuV0VkXX2ramadrcEE96yinvugMpOqws3NkSgd4Tw54JJ1PO
GENARh5YndAKPQB4GNqHPf/z3CmVe3SVF1piPHlUBO4YK3KkeJQsTeVNhKR4ryhkyqtYcGAnzdPJ
m3Big+mIQHCTQS5YtOgniypufdlFLjIXOBWZHY+A+o6tt6nrJFhX4hxFA6qI+SC1yniX0cRkpV1c
ywHvvmZ4DpIFZUKl7h303+gazGQJUKnt07z0n1icJQdlM6+pt5XciPjw1/g4z8QUyww2/5Ba+ssy
XKUu86bcVjOF8dmtDAo8l6pMDoJXavTStbMSgyqudFRGfmJiZClIfQJ2eFtbRyjk+xVN0xRu5mCZ
s/nj28yqQ5GW/KE9BIq2NWbh4DM63CSgHVGE3dkbYL6DRDxGYltJbLd2Kn7GhZ/syDmCD0+NjJgV
xKHOi8wpMhtdxxjFARoGfLYhW/45NVB+4OD1YXHv0cO/Df7BsuSxxZr2ZT8Yipk/e16sq1triBI4
0+LW47S91pvDrxIQwIR2Qr8Njnmdhak4DPHWDFqurYMs8unFxQUGYFu1H4+oC2BjAVdnUDUmBssO
xv+ih+9oJhEPH+dPL6sR8TjxtrEVzS88+fp8NeANdOqSN66jrRM8xoEdcFY9u5psPVLVllWXdtJ0
ACuMr8A0Wqsul20JerOhx1M3Pbn+T1z7fUaHrIesEwAaMaDV2IWANb9bnlVD8h1MwFyLUkZEZXDS
2CSowo1j9dNfLgI2zfiHOvhuFollOUFP6Ct6qTnxD4dMYVz4oYqE9yM/+Uvd7WDIS3qjl0mczV7h
Cv1RuF9/ZJNHltCGYMtmP/vhMURBC0+2ecHoSlfKMqnkLZ7RwOOStpb0XEl848YZ/j2uvAsCSVVP
8d0FpRf64nAFmAMVmNJ27+LwlOzlqbQiV8meJbrH9Ud1JiAOc8DYBw4K5xCGHOVcwVrXShrZVrwK
2M8hGqlhcN/xU1WUYJcaesTWDAuImI0dS+tFIwssSAOiVo2RtQXFmB0BUTuF/xvPVfE53R6TAkWX
FILOt+4EC7Bb9pcZBni587KCH99eHlVV+rWG8j97OOlp3hSWKzITOlPUSW/ER53fDSoBY8k7Fvpy
BI/r4bGtxn07ppzNjfwpgwpwssHiPorSgF2tr/ygqlBsMDXRC2Pqghed/ekwDvaQUGBmFTRb5r1D
Ki5hLpAZL8YNmfgOth5kj9tNNKH6tKz4VFVdWxiapYn5b5giNekbmMUFCEH77MUNvMaQXD0JSq+R
7OV0O4LKkQKO+ihvKS6GUHVoBbx2ileUqT+vNbVCKYxz4db/kHwrMVXQ3cf7oeyiECfCiABpr1ZM
ytb+Fk3NXv64B5Lv93aT2bUoT436QO5sVRVQrsStZQV945ArIrL44C7JgWOUTW8ExHIBaB9bhh6s
iK+PSPeBKeOuYYm55UcT83kuooc7nerxBzzCaJylbyGEbZ2bF1e0lXfqO1PXhOP8D2czQzp7koDN
hjRAisFOkUKkdnJ1xvJ6JeeTFTYy1d0358hss0K/0uJxi4mQxnLbUhMk2RNNe5N1iDew/7QWzUwd
s0ZfF8A8y63Jld9n93+TNhZdp7EekIZClfgQIxxXPFRVQQn9h9P7fjMeoj7Qs1sNbhRD3PfoqxiZ
xilY9ktZ4tw36U7WIzjCvkGYWhFYroLS0wSltr8wHEnnykUtTeG38fM7Xzb4zocieBmmIuR0CDF4
NBa3VczLRZSze7PQe7iQziW1oFg8suvcV3xqdiOLd8bGgRjvZ5Un8808uNXz7M5DvOf7gGPl33Rx
P86C5FSfel4/LXEOEpx3FX16i21FEy2uwa08L7KzeVsQ3SbPqoTRX79qBXO8cer55nZHVBr7lC99
Q5XOP0jSTot975rsfTW1MvVUNwXlJkKryjalIFXhc1jxcYc6DnY8Es4CbO8btmuudZvWrSwwLI3H
Mz5BK4xhpgQqCKoEP8pKpmAC56DRZO3Taji0lpHK9DUZ52uFsu0+FqKOM4MsSNR4KD5yOz3IJzKR
nBZl9+ZTyqXtqoVtKq8Nh94e+vVPFZuc6a8EGirCoEFzCurKuJefWqewtVknvNOhbakfvitz43DQ
qID1zyLV2nrCvz4UF021ROHhCPVChFtA2dDFPqBbyHZdUoVRHFbR5utF2QF0/+Alqj/4aGiHDQeY
XjJDSVusiDTaeew0WOi08hcTpdZJE+275TSO29dJOXYQb4SIVJMJ3Ug2XyU5d4HvshLWZjAVdxEa
DwNZFJyTH9d9yFG7HehvPbq5Ymxcfimorcdkv8WaAuIUtjSIGfFmEkZdopVVRrnie54OtNJ+EGVz
s9MDHL9H7+teobfCt2zCVjrs+/WvdB3tUo7ZPE/VOrcZH+iZ1JkCkmlVVngcVcHqLMGEv9AOpXPO
pLohVZcWEC8pfgtt+meCt+uo6gD3vmeZupM0K+nflzkGujOPDBIQnY/CjABLxdF2gfZVOW5f1GbK
aeADju5WhovTOW2PyP+X/4xF+N7EYVQpComhqEbR3UlKwMb12t8f3puKC+16hoWw/l+9xpQrFXJz
J0RBw+CziUcc2WHYrf3EAUZgHSJB5M/oF5ou92kR1ec7yrqVBiPYyjXaJXQzi5onR7sPxPqItyun
coQwzn5IaMiDhnWrWUs4ZU0Y4QybWKCnjFPa9ctu6QXbfjMZYgrhDuxnLAV8Kkc2dJg29IC0gKWF
jv+LtT85Hf7hEuo0fMfaCzvksfTXzmQOGnxdYcvlmtdqO4PQrgP+lN1Wynq53DuB48IEr1xaKBRo
RAjofGARv3htU0vhrw1H/bf9MRFCEezYwZI5j9x/tcvofFuLfgJAixDmZlsQwPCeuA7WwUO9n7Fv
/6PYzUNTBvs5GwQ/0AbZJNBP7XrL3+YaB5P+68KymlrtMpvYF+7lkGw8kqZPyMW6iBWSd3UsVm0Y
ZihR1hkeAocEs+Yp9RcoHkZt6mreJvbpJ2MgBMz2mHuuH75aTsTzNQ7rvQVhqP5BCfvD0eLwEaUm
ZDd2HyDJcpqpshs7LzRBb2i1XuLWt6CGi6g2IaRaZjT1NcUju5aTHFDXRv/nO3obIZxvJkV4lttK
qIKIWh7qd1wJsQyHiAxs1AUEt4de6bbBr/E1Sh/LcJSE/coEtewJK/ASei7nxg2kD8P0qlf/970a
l99MEfQHhxgMAtsDutSXc8KQZP+pa4jHmH7xmuDJm+pWBv3dwZeizQi4d3TnaG7O/Xr4zGDqzOjl
fr0SC07vSpjOa9G9qe9r8gwZbhKKS//CcXPzxcb9r/hItF3Sbjv2m6aB1Gee+Znz15fLXYo4yoVE
Dr0+pYLNBZ384iUH+QP8NOJ3TdV2z4KTX8lhfAyiK0dPLj22pR78p8PIU14KXf2wxyHzVgqltSrv
XmhgO28eLgr91MWp+kR2V/URDjLnGyaWhadJyWnt+W3rFsYVuG7+PqH+OtHizkGcTS8hNeMXvGLi
35HtycjHXkjAuwOucgSe46u9MtkrRdU9v+gPZnS/ntTFfvo5fO1U5/TodTeEG+q5drPJ+EeY1LTF
ATR3rI0B8bDQuSQbL0vqez2b79Z3OvVr5+B9ur5a+WtCtDU19uFkBLU334uCJtKyClhfm2wqk9fN
oRyo9Exnro9Knb5Er6o5V9UN4WzCyG/K3vXY+KOhQLQvuUuCPyFfn41RakaoEdQNcMx/lBEiBH3j
y2LeFJSvSqonPyJTE3ee7i/f0R0IemO3Y6QZw9NzJNyfTl3OQWZWiOMWUT83ZaTpnxbQoRxMlOn7
1bZthUVQ09zk7hDwz6n8sm2GbRICU1PB+QQ57WJzII/UvJ5sasv9FFp5NaoE2yN3uR3bCXR1Zj9R
t6XBH52wbIoZzbUF4SnFOWOiQ82LOjg0S/mBYEGtyOoxOebTirT+y8l9LV00gu9hsKBz5nvVxLMN
P/U+7cbAKKhB63fUh8yQlAtufqe/cqr47xefdLIHGPn6rsQY+ShKIFgt7ZE8ljyAKGQP3gGSYCDQ
lkdoUSeGuCTuQBXrJ/c09yjWb5xh9nJ36fNEocPOcPE95GfSJp9qmiFazWGuFZ8ByqThL9T0SBMH
5tF8h7B4HPGit3VEaEpLJxGmL9GIYt/EO320bm9KRjzx3uMh33huEodpQ6fY0EaM180VC8KrCb2B
M5kouk+g0viRyD0Wq8UAgjMEcL8EHPbUBpxgYEy25OASg0OTIWE6ebQR4xKBhHRCfHwgG7xP4CfH
xJfZrqaWxlo8Gu5ncB+OAabesUrrtty2oj1+nlOCctl8pWYJezcrVtMPrs6n2sSRy4ujq6f/r+Jk
FwDmT51tYApilr61XfdyytdlOUSv6okJtHTWUVXMqW4pRqkqEmeJ06WZ63JqDF2xz9DR4IxxxtMl
HYJintMHUtyzClax8p7NEyVlK8Yfjajp2JW5Lc4Uj7JCSYv/IVP1ZW8b6PWton/vMqr9TIP19jVc
PyPmRDO3kgEV00lOGY8Ub8K6s1pGgKgC7TYtchtDElA6TSwUvzgLfyyVw2UteOQlOIkrTZL8JIha
dMf4lZRV63Qfso9awuL2Stg4ITz46qcg9fweNg/9jcHGzNfb6NXqeVGREk7jldfMY/cDNN6CCLKG
PCRs8OOrAlgcGnEyOzKVE3e1B5i5uEraIDOEqQVywLd/8CYd5325hsgY3EH5XGkJlMA1A9vBnkKR
rxm3OyvxnaSel+KpU/frZmcLAaqROLh83MEzEG0E67F0WY3+KtS6Y+8x7S2gJKTHRZGDrYMBQ5/p
wi6VS0kEC39Y9Sq2r5v/02cNzGT1TcBSwR9MhMmthkHKW1Rt6ZsPVcwin7fxEItFDLNUr9PrCqK+
1EdfwKk3V1aVlY6vdRHwqlRfwJ1gwXh3EYD5Cyxd0JKjn8thnh3P08eJ+wtUp9vN1ldXN/HKBMIf
DfjWjOP/gwsopK9urkdRyRYJVO1sXuC9ToLVcb8K1oVTUzNiulesAjPzpD5roaLUtK06mw3M10fB
87o05o768qrKTVYx2NNtV6hErwMQl5tpia0GBPhKQHVb2e2dYMnVvQXM1Z+6sjiizTs3Mjp08UvQ
FZMKviXbaizFQpeqeNfN5IRVMytR8I5xuU9/5FyKLRKz5R7gU3/D4nvMeTzl3mHkRwNF2vSo/xEk
etEB9DNg/xIqAWkiaX/0zNlo6A+aWDz4Hi6m1fkJaczoZqYeywjrAuIhpN8iiv5i8ZtGOFEBrTtb
c1FzfFzUCSD5mQjhfVMvLNFeh5eje4OMZl4ZcslCqDQPheK6Y3JH1WcGnGXM1QMWLA/X0djeGd5i
ys1WeIC4xrLm/nwwFmr+Czse6x/XmH7LULVkxRnTliwYHc0L16KCbgi84Oes9EvZ2HIca9gKs6ft
O9RpKTsrh9ixghiyLbvpQ6DWYLxfeq/pFCl6BWNA8upEtr0IDeot9XEtAzHiL+fq/Igx6c+OfsPI
QtNPGafqeDVpxtU9mZJ2y7FK4FPJ5oSYSu33RHuKYEHMQoKoB5mg7OM7fdXyHMf1oskgdUkhrS5+
E6HXw/QrYm783YnMsbzo3gY78KvI1mzlcsqnHj2BQODnShaBQrtumFYxqsWlimykNaxh9n6/BKND
zazXkrcApx8pqEc3AFm74DiFkzDXdeHS7zE7X6Jh6TJPIrreMs+0PlyG3hpaJIJAmty5M/7sVyD7
IpVGDLU2rncBk104zIk/KF6SGnDbfsMI8Idl66awAZBZdlHIwFrsiF7DoS5ZFr/iknUMAG6JtbjA
/FGOBQ65aHfSCaak1BG8+ubk/UVyIt2cEkZyfd57wQEtm3hBV2QxJQqcBARDJF6uSra2vK1J+mj5
B1ug9QLch79BT412Dq55ZgaOSMYXegLcmC9nX7ba1E6DEejRZXcYZTQQmffsDplYeOO86OJ32CHJ
G5qOYeq00nYcGtU5Wq7nmEbFiNT/y6nOZQ7OG0Hy7Gfm3hAVZx3OradiSStXcnkhjGv+Xi0E+4St
+Gi9Oc+BYGhbl1xM4z8k3xVPRPwXUPMDn5eYm1lqqomcTfRMajLymGHuUjDnxIaEMn+fmaPbC84E
BvcVTI9c7zj3mpD+4UlB2tEitT8GbBWn6j/EZ/IX1wmAumJFSgAW5mqntCzMKyjZiPD8gHIMXrhH
wkEBktj/QQpxX183EiGVxncxYI9QmfD4EgB35lZCq6SfHPoc+YGPVc70w7QIH796bQ1o8MkXvwYP
jxo4dFpVl8xksc6NS18ntwg0NDfbBFwFCCtRlc4TAEhY2MTTYb9DDx0m9g0G7mcKkaHhYD+yB15V
9JGO725S5sP/P9uwbyqI6kQq6lYLu24VpVbZsIVQTcab+yQ5tgrGt5/CzbnH+wktMipSOuV+QCiI
3RxxPU4X7r6IEv7P9ARQcRuW2/7PaecoeL/GMs2orxz18vI9UIqM3dixIdq0cvxWzeQpL74roghV
QAw05REk0VedJ4zR4fVLW0waEP0izoxw9+obUFvzGCe2JfFU7FVb1ICdAFJ4v+gLFrKnx4c4CuMy
cizGZXG4eTo3XJFqRWGoF48gEqtQJuxOkBWz6i7wiXdGEQ4o4gDxVQxV2ARXRVRPis1RXrYCzc9b
4Om1DAXG8p0OQnIS+nAjcA1n7U3wwm24cR1oRY7vBF+nQaQwvu3pjzFOHnr+ljEkpAoL6MTSPUBQ
zBi+zU3q7bt2oE0LgdJEaER15Z3Px8EL0VQ7LWLUa9wLQr3JHieoiRzzj3XjB4Cn5Gte9w+dSA+L
liRvxODnRwZQN5SUgimQkfpBElYZ7/6AO2oXzkMFg3p9MSR/bqX+YIBtPHfUYjpCTKMD2+D/U9gE
WiRtw+EHwxUyCBTWKjbMxxxcMrJWje+oxtPgb/U5Wu59lYfd+NNSz3VDAKzGZFD996fX8AW/L0Su
2pP/Iiv9//aTFnOV0APX4YfjmL3oDtXfhA8F7HgB9VXLtpj0oOUIQeclF2Tdqojjl7OyFYzFGt52
xy74SMpZPFJyBW8eevdVDW2dajCiw+O82crG8htSQv3l4Ia94S5hi8SiT0HI3/WAhkpxWbizrF5X
NYw42iXGRxdMoFeko65M1CI7D0kAlWTdNcD6j9PHbpUH8/FsgCqYSlm0yfUzYTkoiVi2fKo+8U7S
y08W3a1Sxg3j2LKSx4zypB+QK7pq2G3St9dLBeoOs1hNf0nrP8ckuw7UhxmOfhu85RkxaNffku12
49lEUIuyw0nxGJzsVYS2QLhiWveVw636vXfa5SMtVh1n2bO0WX8Vf5GlgtL1c+ecu4457V0n8Q/t
3pAGTUBeqcdCZylJNmHeFCf7uigzSO63h5UuHbUSiWuTjl6ZxMTee1FU2bPc8FFR8UCJ4mJxT4KL
s1vZE5vljTLsmL7ZSXgvPsBKEnXFbFG7M5g90RcYwgcO9edMah/UBvY3R8vC3Bigt3yLIb4n/YXw
F+s3ZhtSfPar0VVjmDU3wu+382OEwt3PueNPTtw0JaLHViASSmkE+uWr4AfIjzLxUaPnEuccviia
7GLs4wEPnTa2OEqlNEiGbtxAS4iDXHKS9GDkFXDKC7vP7C+8L0JDcPxc6kWo+ZeseEEg/uf/8/Xp
uVEcWNmoS8Vqp1fEYAfS4yRIG/hhDitcUJJF37Ci8dTHI1ofmYN7K/6mAqY3UUYj67TagRz6WdSE
juRIUn4wc7cLhhILMm92pBWxPR+iTwOdG6Momy9E5uW1Xw0PHDdtDDL/+YqQpJ3y+C6P+mvdz//u
0SzjJjGjnOCFjDPUCYWsY8+yCPY4fdSva74eESj1EQfO4O1OEgWFD0Q0tyEKsraJc6/UxHLcKBFr
VMnVLoRt6kPNcovdMo7AkxI85HKYSLU1xIiD0sO0HX+e4wD/jXPdDj6R7OwIrJPTO4dnZf3CP3xZ
X6UNG0XeG1sus2UQUwqDfltxIJ43tz8FLdE4HzBtH4ZUigr5bjtJP2TW/PzlQcoL+kHImmLmByYq
qCq/zGs/2lWAiosyOeehJh3PQlgiG38DLFkYPEGGg05d13shA52tqdV1LCXCxSMZO4Kw7BFzzgjr
yvoExuYWgSjPeCntn80CpwS4WY3cFRicRN3AXJYSglH6KwfHnRFb77+bCPQ7EB+f1kZKbnKC7jjr
jowtgesxicFyBXXvJunx+vHODfhkHih/yjpL8AC4OPwWUsMjen3zBwy3/PDCMb2uSPf6cFIQ1g3i
7jiBd9pDxV022XIy8Ok1waZFVo9BKSMf9wW7c1rYkMFA/qxgWpnun2YfAAac6zS31jgFFfnzV1/F
iDAG4Dysdmit7SDQ79Bvk5y6cO7e3wpZTuN/9YkVh3cQaj0R0lBfQVIpRSW6AWAKFmicWR50n769
+cLz0VFq27XLJWNOLlsma6ptQAx65d1h+PxqIAFXMWfRcyM5kMNpchsVl2Ja5p/x9x+21fufZ4YH
KFqk3IksZNJ0YgsCp5g2Mti2aNrSDtp6sQS9QS0R5rXkFEpaTFPZrHiL0wWezakUKSvVcL4bWSHD
OtnpvzjyJZEjkp9VKkvABHJWr0GAkY6QZJeaH9IvGaY+C981dyCM9zsq8iI0+rI0sZ15M7VCaKHc
pCSKvYyUzRIRqy+gyUgojlEQYQH+GtYohsDN337U39z7LAjPK76C/+3s6rV+MgW9QkiD3+ZM2vOl
kLKc/Uz7JZuiNCp9tfH7AO9Y63twcoTsNT5H4PHuzivNLKxvUJqmC6yiJYAICLv+u8r0XFntIwDl
sW7S1QYtIplWgsG94Lz5uZTeNjEU58W+0sYG2uW8TIV+9Oy7mJpKjBcA3KHdNpb2IfJAS2mRlETk
5UYCVOGr+i4wtPEXAivfSBIXGHaGqi1E8mQPYo47+GRuXMbNRsOC9Idwoy92E90GHCScDICNa9RE
zXPhqqPVZQTzRkDqDQ6pxUgYA+pgBgvH7f11IVqTxav3vc2+i7w+0hj1BVboH7nRd+L/qAZd1HLP
xwET1tbmqzSmU+uNfmwFVa+QOfCTKEb21j78B7083wjnA3gqNvdUDsjJfAV646Q4vgpn66HcRtmO
KtWU82fXxY1EWn3khPpdTfLWn3LUl2g9+hBb4pNyHMpHhV5lqjPFcCiV9pLx9FZ9AAmq/z/steVP
jnIgvVZh7ZjXyCDQyvJVQzFpg20GVu6h5056PiMXmnhqntk+EYuy0jH22tr6fhhtylAFTyUJDDri
8oGY+qupASwl0s2SQVBQ257Ct6z7pzdcs1zwmUFyLeigglCkuhZFtCQOj4c4+FlxA+QmDt8rJeyf
UQJptOIaOop0n1UvQWHm/afX0cCR42JmLJaKq6yjY9loW9a/sdFJMofctFRSA+zC5RecQghbWk/1
KTAh5WdwH7ifsj/qYnXrlWh17C5kRs8w3KwFLSMLvTJPaUrUVfUI/MNLXAxlehZrSEPLn6i1isfP
wd6btGV+osZnKg5rIWNaq7Sqxk7oKAN2Xzfev+jqaoDP0LlCXF9+38UdacBX9vXTVrguJL4QGFFT
RHj/YU+RvAp/LtTXrGJ43vkCIeGv9kn6R/T1Cmxa1DsEEDGulg1GTpmVEXsUJCX9xXdyHPxZycgl
4UBBVZTH6j9ISVfkv2fjEE7GWDcKvYWjj7lDbqDr1fNCJKqUqRG8UWAwTbyOvBF83VflAQ1A8d5/
KHI+DF7wvchgj5PxdB9jfH16csLF7z5cDu2EcjuVFpvt2QVZAZPG/WGphNVve4TSWNQhuTWijlsS
c/wVCbMuo5jg6pRvRfMpd3u1v2O32irvE7RO+s0wkfQCWrTNQEAMbXrzj4V5UyLERAcrv3v/BpSS
Uh97aiDjLkwK/rz7LC5ipsVtUgLhLStsfVDE7VQVbkuhTwlpnXKWH1mwBgVnaFOnOobnIOcwkU3U
+kIvvu9Og3CXcwE/X8aMK8CGOVGWRtktYj8mm92zpfg0l9sEpWclaWms8I2sfoPBNvMCOQWzvg1Q
2efnH6x5kxTY5bjjGboXFBquMfscxZEh2Upiwc+ZQ1lGTHHrBhilZoWnfeGio5ftr2bWaqVj/p1+
6ByMfS4HagQ4C5er7Gnuo3zuUq3cEz5YGjOinEq61I+I5fZncs0D595rzp9VC9V1gE1Ik8wrhRtn
MBjXnmJQooMBuEJZdChIjJjJ36X/s+pIbdCJnrHd2VQ4UMjxRP+KvsFt72VoV4oVRGh8wuSxF5uI
wbdbnCZkWXRNFvSbOoWbJddD31fhbJs2R0JrJyGCDaiVJk4Vs3xxt+kORmqhRrrZArehX6Sp9q8h
VjMyPRIUqNZxJQjGRWTlB8iOF2yq04byF/PkhkE4xEbEQl9zwgh1VbwhGWY/ryoTGny+gU++NVda
QS3rcKnXbm00oemBL6qTeYcM7KgFXFHJBt00dFczfSC+yY4wtFe7dtT+yuXe7jsca7s8RHjqeM5R
Y6unsLeZg07ydxvV4MKypii1Ygs889sSEZwK08D60X5RvY2atefAT2jWZJGAFyufhPkeDNi3bU0w
4DvxQlGzO8n9HJmk/MdbUSXZMlwREnHlb5BWMZQXAkaWp5pFujnkXiBPwn2NRpNsWwvuDzwnyRi+
JSq2/FGnWTrj4i5RlVPG1c7xHAdngLGKxlENpdru4u8wyQ7Euvp2//dgFeex42Kc8SuBjIYGLqcG
MD5VWpdXjVsyJTGHxKD6LoKXOoG/NlI3XbOFrk6e+R7zl8q4kk6aryX7wyFaJWrCpZuGQ7JpRUSm
2vwqA0YUtBqC9Pg0/0Rhz/kkYV9aRwzLQUgsxBGb1ysOMg9S3rmep1HD97UDDw3xRq0uqu7haKHL
qgrieO2tGKNkex3kU7lxufusC7uIvSoK4hTw46JV0EPHs1WGeipiNQN7Bfdte2wB6QYYILz6MKcw
hg1Vca7xdvRtDCSJkVGgiH8RMxhv3RJs1uLtoQSS9IArpC11TtlMFeDc8xUZJULx1Pw1ycbmvrlA
mS3twwIjnmDrWn2E+nl94IadkTDWOxVUlQWc6tkTVB+7xb0mX6Av8+aV4gYAsSw3qnvRf01N4lp1
8LMTWlgK1oO2m5jWenaEIpZpqsAaN5OeCNPXpP0J34Lm9M7pbKugVsQ/xc5Vzl9FkRmZpz2sqXrv
NaMBtURWG2gphzsj/2zUt/z3YnNkirjCjUTUYCSzDXDfZIsl0vfjdWhPdRcKwRL0dhfqKlBfXd7u
+0Lvdu2QAU9iLBNyT9YcqiB9YvgjD920l9U72P+Tscst19raKoQgBEc7SmzIQhmCoz91FCWs3axr
K5pNwcTYRGXyFmIcm56fdiMDDGDzRuFAMhbltohHL5QzHTJCUFO0aE1pNV+kuHZ5XgnjKCLTbhzE
MO9eINk8/4THMEGWFlgkb+EHUY+QNoiqSP56RvUB9qhlxUMg8id716IMyMr3KIZGEqd4fd8cTt9a
SV4W5V/anWz0027/Cu3bw1qq10r7htfVzJy+U3LNemSWfHn7QzQXeH+AqOibBlpiYyd+0ktoClEo
ZgEykXCxp+KIkg8RNRnHIK9/8sII/ZfE7r+TXEw5BvPLgzorFzm5p7NCRLtWmt6Z8iO76vHkr0kJ
93xxyG4dqG5zSWVnU8o3b9lYxReySbuO/fbmBEbcCqmLprZnuhCadUuvG12zouHJ+JXlCIUfbd4m
47e+b/hv7JNIXPz40Qug81wfJ5iVooBJG9hat7egkz+HvTHnHsvCxVXz6DoM9qfigpercni8rOe4
u4qQ/CcP8KL3iRHVDaoa1E+ShveBpIQuXOSjINXsvlup+VU4R0wFyuVVWb2n/F0pDhe3AyRBvAoa
ZWCy3uyVPlyW6UIs4KodJCBq6a/gUf54YdLGC22+1HJtK7RAuUTBvbfmF50os4hoP3mFX86KiTgQ
cidLErmlxuq9P7V4deAB9jpdevAKSPLim2BhdUFwgS+6dHP45ych93AE16iXooApr9DEqPaZskpx
e07a8Z3VDgCBYtvR5PMSkrihhRz4MQLWZDCMqt43EyaYbcULmDFonPpDQ5oVBAEouyrT3/Q2Yjs7
zUZwM+cSEHcD5XJiDUur41iQYwzxQ408bfxZlbVAOZyhwbjkaBjSlP/bJuscV/l5mCE7KcOI7M5c
QCf0P+B4I3HT5bMnwRcXhW2YtJkMLiNCXXTI/agVJN+HB7s+gQjuh6xGdNZFA7T5OBabB7moPqyg
Cfi3rsSl1Ojt259iXWizafBqO9KYUrkroaoCHOCgMWISnYq2EBNDVdHK88mmF72uLe0UriE/8u0J
la+Nf7kAJkvrlCP75/nWynFsMa6jQxv4/SOOeC66BvrebJrCy8c2Wt9htx1ZNdV38ooFNK7AC/uc
H7kAnHq4xwx0WaopbW7eYI/VK1+Ee/5oVA6uWZwEKGTPkrX7e4pE2MnBMdU4iC+e1lNNrTOi0HJi
AV2x9l5tJ6eIr6Xy+Gj5T32JLzIPcevIOsCmGhwC4oCEGcsVbwRkpTEoOrMVd9XR6iNRxss/jghI
8hVEPF8N/4XzCi+Z/eBtUu7dxBiwmcVBt+Q/rLErbMe2H9zTZhX5jFELZ97bdX81xc5c/umR6L/z
RhoK1bT62us2XJeZn0O3prWJF8Hk4q3G1vHB5bLWJwsqHAyIVTiDGyRIEvINrKkdCgpJffiWxJG1
539RfQuCAFLkUpWGFKigPu9EDl3xSAvTkiI+cPXQ5rEf8cCEfYdNi5spfHrTHJs+mjXH7qTQU08/
xRox3QycuJUmgKeujemzBtXY7rxFd5etFOW8upoYNS0bKN/zXw8VlPDW6H1Zb7oSddTWedLrXhFO
S7ANoPJcCD+k6Pu0glE+82EVGJWfxJ0auQm/E/YctB1bI/bzcSq5oajhkneAgKo2Ere0mUuqv/eg
VSXNwBjNuRmtP+5FZWqrH46Ru6KVXKMjCzh/V8FvmaNkdUoBBxFzjhQNvrF69KylhEQt0WuuJOy5
6Z2NBkzMkwLKhA4chqsj9nLpWcWSZpfAwSz21xF9okn1XK88B1LkRCuTy1jMqK2vzTMoM8V7/qjL
wHv8DEOI3l71uRJdH5Yb+sZKbvQQRJcp2FPGnnS3cc27ErB1ctREUlqC1CQ0eIrkADOZwlw2IAcx
qbbi9/r66U37HvMj92aOxD68yQhkpAYxfX2Wrtf5Q4/ZWxrnROCwLGWY4quU/8YvEFwZb4N7v8C+
D+3AFeohUZwMX9He0S8x9BpCeW4Ttjq6QOYU18OFcvk3a8hnvJfGNgG51rIj+05TJVoYVEobW4M1
4U6yKzngyZ7+31FG3GPEtTWOw/PaMFppVUSUGdOietVMNL7qMdhOT3rWWYLWxYvgPTChPvy3o2/y
THl2fKe54MiO+0Fx+45heZ8kSFn3bbBU+UFA76p4laysnLn21NXSxTJ59/WwQcgwWtMvXNzQTPMV
AI6IbMAcOPIHIhKxr1LXFyD+UQusJ3iSa6a9spE3pQNTY7ZxL7AcMztkBRcbRVGblGeMmopKgFQm
Pe5mAQVBd0eb1KjCmljt+sYcPT3N0gBvhKnK3/ML0lV4i6Di8VUl2C0IOk5Sdxs/xWQdOsneNn5S
JR7vy/0eMEkO7TJ5f5+j9ncAS4MlsQmtuyPvRsptzg26Ev06NMe4Nwh8u5o51j03iehmM77QbUgp
barL9y6NpzzRGPZsa1+9tj64EyZf3YJvG/eBg3N8yg20bdhZ1VRH0Uo5s3cy/IdVKG3iVjWt4dAK
j/ax88QD3Rrv+TN7q6GAOGKdr2cFQo2prssmIFL/nxPbpfKdKtCl80plhEY4vn+vjSJM+toq70St
/dV+ecCMNkmZBCNeJrz225u47Iv9Gi6UYyhTw+n2saZKbwUTpToUL6np73rVpAttPiB+2BPUtYnc
vLJXXBdKYmSucliYPmwY+0Hci3eaY/BwpMvnIj+Yj/XjPvz8gWn7k7i43sOHxvGVepwQl9nkeQmz
BNxMOMW0GljbIFhT19LGVc5vdjUBCqMwYT/nEJCjOlI1lx1pWan1+nQqmdzBpTOgjxViTi+x7+VR
lGmrUaWEV2C+OFbUue83rHAN8rTNe13ubWdCBKpaREE+Bdl7Yn8K/wTjAsLxkRmcQptBwLb4e+Va
e/slYRj/kV+Qumr2EstlUf0sqDN+SCFbbcLnhC1PgG25ktttksJhgWhBM4e31K1H91NqA1HD1oF4
nlPdPjzfLtYI01iXxRmOVAYJLS94aa5+SDQTAT4mCP7ZQHtcJcka3eKiFfiCndDqyQiviYrVWfT8
WElp0Xy3dFwpxKDYIQvhE6OIjfAsmGMROExoLnoV3TCsnNmwRVXHNsTva8/LO4rILw+TlYrK9Zw+
/P0keXIUF7Mi9EDyrZOmI/9M33Jx6hsOjo6mtKEem9xTwdX5LR82yj71KcN8DJ1LpKjCzZEU4OIJ
x4HJGa457nDaDD5e/YZxC4smC4zc5CU9HC77cfB7ElntZ7JetVYGJm7PsJqSYTozQYIH+FrMX5fN
gUREXOj2N+VnIZdwCwOErMEpJRFRh2RPe+770qLyGXe7RsoygnQRHJm7R26m49w51UD6jWaD8dco
kQCup6gJiY48DmVWa/II8wVY94pB58ITcRLLkCpfiddVo54tbXuCM+WBFeIL9XUyonU8xthQ7aBA
RarKXSK0rDt43Ff2E/0LyC2tU7QLk94u9ybcDo4vHYpIYAyeXwAE2o6vcnzVjWVgslXORiEGqBvo
1/xVS7h0fxgtEj2fc41o3ima1KV4EotqBCT+alfkoPm1aC6dBYLd0E/sC0UcJY6NyB9GjCPpXSLK
L2XRcBPfFK0GqdD/SYG9W4VrFtwD6LLxIEnsD4flqtxxfb+My9f0drIIPSGfZ+DmlD9wC7itDSNg
VK7uyAsprddu/cYKFvMNXd3ZqJ76qrplJzzyf1aQfx9u9AHXCAso3dmZCRvkqvFR1wPWGkCCSoOt
XdPHqYvQ7mIEvQEKxI3IPoDiFuXqNiyf/5ELFDRUO7UBTssAzhdXoacnlEohtx474rJYqbrGXds5
z9zT12Sciho5ua0XhRZEeznBDfsB0r9qghmNluHfyAAqq2f/0Mq608p9B93n+QW8IgiDUa1qqa++
Gjdmjhe339rzwESQ3cUGeZiCODt5URaGgMX2Whx6h9xq6I5FCgx58MFblC5IG7Nwfbz+mcC+eH+o
WFHZrIAbtTrgqI3AOgmjm26ntge/+zVMk2U9qT4wvKp5tNLGKgq3ZiOmaaraVWS8DCT9uodl5KCQ
hycAwD4nC5VFO8iMEutaKh+hqm1QhwkY34vIb2ZvJ9vyoOWmm0M9AEdCpZukZTLg+9E3iOjeMinD
7yMiikzDXS4Tgd9sPuCMDftvwubcKLz7wAau1HPz52+NO+CjOWjzVx9skuur/UFXJ/4CKnYsVrZU
YMj5HSPaANa+BpWpEx7VjlshCrrg+GriHhtAb2goSn1GPeYPExFCT+Mp93FgS82bLU0tWRsHw/74
Bt2hsyGWcVr4ccltkWO0UA5eiZZVVgDxSGKNyYZ1XWH1yKQ+GV2G1Ptv6xXqjEQFLFDXSvmb9Asw
2lG02D4eb5sFETQ9unN4YyOiJO+k9zZPnM2AQbyYldjMbF2JjAAoIK2WBw7YUzzQv3AUjwkAigHu
YyIGa9j9P/Y8lQmRMeT2+QwGbT7NIKsH4SvnfGccPFAVOBgT43HyQ2BlAraDro4mMv0kn6oadHb3
PeKXbNU13CWLVc9PbL2Mjk3FAQ69AQpuTy/rWKn0mngBEtIHgE772gtzInicnaKwzFAN3bXxf1E4
HZuHhKoXmn5uTWb/zoS1Bsw21l8ImiGUzDJHYnvETgfY7K6pUG3LdjmFFCqaIRrvvKxmYtVbwizs
b6UBDodtuQEwCm9vbjLY4I6DK43NICBJznWPTaSKJoK51k8I6hyGxr1T87xYW4wCzSZmx7ntfYg6
Ev/OGxs2nOHZTLliwJ68TTwE/0edZAO9/bQJCW25JcnzlF0yNuSvgeeAWXJJCtj7EJnUkcRcJXmc
6k9BTljiEC133FJX6QGFnh4aasND2phdH995sre5AWIg8iDjdu6ODCea8B29nabS5gPZ6s+61DEg
d1BNApSDaFkx+9h7VhbKJ3szVNEwGQJxTvtjDua0cb+Kg0Lvp4Ebg+WHVddJqzu1vMsutk01rMhs
qp+CA8V5GtdpQJSGXwtCIlX3a8hoQ1fMuCjJusRaN3HAucnYN/H3C/0DZUu4v3/9EIU/V5Oknl0K
WR8IcHvgtj1Ji0nvJiVRG4c9MqXejumQTp+rb/IpwXINiHxE3IZsTCqkI6y1DuEickgggA8F9xfz
1FZr6j52QN7ulMgvDt5Z9OT9JkbTfOg3tvrV8kHZlk5VSqOutWR6LlelHM42XcsOh16vAHaZPprF
X2wlYPD6TVUk9eMNqM+2UaUHZhkp4L3AAWjl2bXkNL6mYWIx1ILhBcs+bGvAexZ5DOGKgDBfkcWf
+mCwf0v5MK9LUPQXZox7hGKzzbz05hgB2uX7eZCKxen4FjPo1wopn123pwwZ821pdEkq3fX0weyA
KUKXhuGBiqgCf7lB6Uiq8+TQqN9CGTE4YauzFZLOIUQ/r0KZBhJ2rzNanWF0Pb4WIxgWYQ4Qe5V3
B+3p7zS5Tk/Zl1In2uUYFg9Q0uo9ag6ap0lLD/J5BS2R5zolsrDqWKzyA+JxQWgCmx/DAyTT4DJP
dBGKRCTZvFhElgm4dWRznEovfwpD2QKNpVO1+VASM90JkB81ePIkczZN9OdewjO6tEMIkZZun/KF
IrvEjzg0AZDuDh8O8l35wnEtccuHwXPNZ3/ImywbuZAnG8tbeCSxsBztNj/0aGrdTh0gNnicbZuY
ITNU0LJinXs3LYzmIWx+cnn0uzMg1hlleuJJt/eYoK4+X6gbOBCa59hXz+bQtSn2Pd0vFxS3CAfR
IgfU48HfCA6QLy2yZBpyzkn3XM9QVvJkBXwEd48HwcJa3w35r5Yrz0Ak2j9aKP59QurPmth7XjGC
b1qwIJ4Bbct1E+yHJm51v+2xJt53oWtgJZqPUILLfFbCS1MxN+7frpT7l3ISZFos9iDLV2JLJ9UF
eqAI2I01Gom4b6Eu4ZZF4PBGD7/ZEPoitb/uHoNNnsriA80tf5zslXcGoJrRtysAszn/7G7HwMgY
ZF1fDyVO2IGpffty9IwLmZZ9EmSSrUXdaymiZNnbVwzNCr/Zgk7ezn0KbUzte3uUYDj/4LktEkvz
jKhidzoA30lfhmgJS+4ojBcygSuPOjZMlVlUgEF3WO9j0Uw0aAdIquVquGqVzz0RAunXItqIOhT6
xo6bdWsfXotXFWRSY+KG2kIn8DI2GY8WaosIxFhqwWv0YtAPaPBi93YU63wVJ1I8+0w0u/rIziXk
gScq3IUCfQvrSFIGXWT9Oa6lhT7dElrvKl1oKaA9j9o5xyoYawE0KVXryDQoNXC5MeI6Knb1AuBp
hkatwLzlAUIUBDg3brQbj60G51AYJ/pos3ltyBVRdrGUOCsELAFg3/w2UHnu4+gYeqp14L5ufpu2
0cO6KYgBLbmtUjRcG2WjjVvQBSReAnGmdwIcQJzhSDMGGH6cYPUCRf2PtHEef1CspKtRqQhQ666e
9F3qE131hFeARI5+cECup8oClRiq0B4U9mSK56n4Bj4BSwskEKhDjR7eD00qJu9qH94W1Ifix+6u
KgaA48F2r9R7kD+YMk0jelfX5dZTH0WEX+rWrPX8fTDkR5spDLNI9wAEZFsUFaDbr8JZBJ5a7pUw
VnkxqTPsfmMtFnC6ziMkpJW+Bsoj0hOBEi505C6sCgJaqt9M+AywJmuRStBJ6ojqhB7FfM+9XK8Z
Fy86bm1PbuORfMzVXMbVmaBcHl5KHpSEfsNFxSDyhf25+SH4jbrJ0ztPdP8SBsGWCAO29Q6E+1Ui
8v3GRM2OZW9DNr5sALiGdd5RUpeUyZ+0OB7bdMBLygXwNdBSVo0OcSo5PT23Odms2RIOp+MnImOU
X12e9TMEOSMj04G5RZyu4wHHqevNzSbHtwJNUszXig8LEGZfyrpbr6029CpPd1LNTK6PvqNVP4MX
DrlQlFuvA6B95re72HQJyxmn8atn2mWPZaGykMIwx+XeUWJCVUkoEJVRJ9LrhJESfcbJn2YLaimc
YsprQRGq8+WFFkshOz23HwLNGIP3CvevUF14m13Ec6r39BSZV6c1m+EXKiLRJyXpzZxQTis5p6rP
gzlC/sQ+w8KjyMbnXN6p+YxkljcLflSbIYsoVrlJTPJ1teocBLSa3nZZDYG3mypntxIeqUPijn99
s+qmMZJfWY29LW91bEKrQv5LBcV7Q0WgjO8s1eJb19MN5QKIQ7hV9qVvlJX28T927O3ZagNyN0wO
oGLGk4gxBtL/UKSX2ZC2HLSdIUrzr9fyge5LVHFuWzlFDNkn1hFxFx6ir7QZ8cjbhlkseb7c1cAE
vvmMeYGs1wyOADxUllpBRykBaywH/x39fd4q2zmlI0rB0sy/HWk+EnKUrpDyK23DHNcXw9v0mES8
kJ6HBxz7LywOXW3aHXZx1ufHFmkABj1Fq1zjOyaXdut83qvETOjUPU3zcXH9o1eGMLo5lSRbXo91
uaCc2I7coSBU26O/ESa6fZuzorltiv4mdE/dMtuY0otTjuSkLfsYdKBjzKOBrxWyKYdJzk8UHpSg
brj6nd3QZxyaDO1v+ZdoLohM9y0awRqULPQl7QFMzcWmRfaplG/RmDb2PE6Fx/DJwXtmLxOLDLEl
ep0s40gVrZ/wC4OBDNexuxuissBK3qmdF4MuN5oo7rcqvvscOdQiawqttIP8ZyYOO11C4A8hlGPV
cT6NPAtaEjHxfJbOj47iXGqHPvgtRwKLyEP4Xezgf7OYUY8X9VgrDhJ/fBMQLyDaKoirR5Zqw5I6
m8qdmL4Y79m8BdaQ2hfDZK6Kt5aQO1wwnGnNMBmWvDLJxkAywW42j0gD5jlKN3EUIK6cEukaf+hW
bEqnOyeOaVucOPh7bGTTdI825olFZRQtKNVlPktnZu5PeL8pBXx192JUgvPVnJDx4N11oKdG/bYI
8mk6YEPEUwPsPbCjkhijhdt/RdYOHmMqa6lwVqRroNFaWGWFKaT5IFdNcXoMmkhHB2oVpmJHbubn
4uGHPEfeHk9VDEbqOcu/K9h1wbhPDYk0Qdn1YYG5wIAf7jbuPh02C7QI/TL37hOud87+QDnNI2W0
eGucKRaBeDafW/Xp6cWXEBQguegcxSbl+R5w34e3yfDyYqJI9b3ySS9ITHeIaUGTbkrivhZQhzYh
Umto+HtuK465w83GSXEk3glH+RY+TnvtdBLkhDjIIOiXvq0xNHVbpnARA+5hgjxCPPCWQqqoWqA0
YfUjcy8fF1xp/IU3z9QsdpOIXrHXNHHQkfWXy0EOe6ZBmtEPASopbxp+ZI+c+CZYhkyHp236GTvP
9O8eurxHwFsMa3CH/6uQMHBqw3wILz9xxhSNC5lHWtlYDOsSC9O13gDkB9fR5ZPYnwnNkjsk06Ve
8fIav547Y1l93hDUb2IGT8BKWxF3/qrzONTVahB39kZLAXeCGJ2/Oow1KM24GIIUBTkGLXDc1Fis
vi+Osc6xDCKnYBYeLe1R5UA7jhCELIVLZFr90BYDeJ7z6lXb0PD2eWf5oX9uDk6H0I6R5Pn4y8Ze
Q/yMl1aYhLM9uTDP0qosD6Nhy3ibbqAxE2Wa3n+1Z+44luiQ40VrBbdl0tYwbHL3oixDr2h8CjEP
cxNaNUxhTEMP/p2NiDuFIo73m2MnkyDaQkz/5TZCsuBOWKsHZPVhd03wdgpU23IEJjley361Z6js
uWRFJmMgdjtxOJhIDOma/Tw5N7hkvYwAgFMIxCztsHZfbdwL9/WdXOKeYHJ4MW9kNarMob6w12s0
kvsVDUY/dWGAzDBfhBELzfbHXzqKBLrKfIfCak4SK8kmHWHTJrGYVlTy1sBbr1Rd6SOz8vt4eqPi
EQVT9vzU3Wyj3NNDdX2Vpkj8WiGjgMf5vTX/QB+YO+KfFxFAlDwIBbTt9cjsdNijTXt+ZF8rJs9f
j9MHh8Xny1jzJ68n1Utb1vrrywB6sfY2owo5IunOTsfWaDlIaKecm77YkGgWtmKFDV2Eu9c9x1YK
Kqc50LsCjgU/q/O3rZ8AcAonfhDoCr/zikS3b7xJowKufxstgWQDMeEfe2qQj0KhjzODGn3AU1kk
u+3FGmpLj6IzxfGAIwkm6D235bxvHRDmTRPsq3bnLqOQNUmSFHa+8syUCoYv3gpz6FsKq+l/2gAj
VA/otyU7pl5dJKCr0p9TmYp9CsgvkO8QBPvX3P1PsuXvS41tgmbsIW4ZcMm5sJLAf/E4uDRKYzi8
exaBICBG6U5/6xi8KKrgM+d8RN3qzBjXtY/PVY2hfmOZToQxCZBlRlpJTkOdn56R5r/LcALlWIeJ
dHwiprqrLLpHKQfVQZOL1AztnCYH4oVzu7fq5kQjmr9sRIcgKd4sifPPdm9s3JDcAG2U7xv5g0op
1WP3P7ouZU2/4FT3UFEuqZX5gvDdDR1oaPNk5z3KBBT/GYy1Ym7jIjvtJO23kBaIxO3Bl8pMcQB3
SBDYRPelY/64LzKFRcZT6TbX2bLMhZuBrzAVgGsquURC6v5jkiIg3p4+AKr5eRnvKpQ0Vnm71+8l
ksmR7WEqEKOKDPXi3uW9eIXXQ5/wPJr7qpjOK2bqQZM3TklxQBokENa41GvFYIA60QRADzrAfgwx
LHN8JqSitNgH241E7TI/ZxFAxB3DJeP15oDSUjo2yZoF+tBKPxG9Ig7TOS3LozFbi5bHXVTnglSd
1LvVFKDoY18lbfPgN5ZvGbnKv9Xa+38ryQNFteAigGWeBhCNzP58EOE/WH3i+Sp+lz1yZxfVXKRb
8N6g4TdGePYItV1pFDKBKZ0lg6m58c+cG/MjnSxM3XL/QP8KsiyXxR4sULKjkdnzjVIwgCkZDjdo
tC2pyueWhePLMBHHvkcF/khogrnmpOdjDW/afbp0oJ9qVLgbkP0qtHbG/oPMmkH7rby7dYhGOZWS
+XFOonn3yqHdoj//ea6TdBVA1evs8m3FTtcxxLbJPP/HB85QHnyA73lbxr7q5Zawb9Rqu3Q0VHj8
zKXfiVJj9ffaJ4MgRpA7l19KDaIsuh2bAH8WgUDrHCu3TY8XXv/ne5ibsZcEsMYRKdJkqFjhruCk
1i45hACTyVth2K0r3lOi5V1v+2PAFR6vUANKwBKOsJ0aXTEvLKNdSa+tRBxZ8kxnlAY5MHmO1FzL
VBrvmG1k3arvjduXGJ97fHBTEg09SG7T8qhfCwvoY0EItON85akd+jZzOEJbBAwjYXK84zzbjVBa
OjlvKv8LDm3cMNvBpgmXU2SAm2rqRipMn8eXR1qwcP8KLcocGwU9C5NPar7/91sS01Ot/uXvgZbr
i02U4uyhy7zCpq2BMDnPnLd6ylRhQdKITAg1D+c+9nrlL+IA0CEQGXjBEOpDdpg1WCTq7YK6LhX/
Gzvr3ykab7vbeNoIfF8XIOo6JbNL5rr+YZwnwylDq+/sBZh2e3TTxfM21EpMZBqE2sk9G2U1Fkmw
6lifNyX/6kE+u1gHMDY1AVqtvrBgQHttGCAWnrLMcxJR+GdF6ZneoYQkstSD7OkGqQkzexwbyC10
5xNBckxoqjk6vpCdDVlsVYT37BRLQzuzI3I7W+x9lUy1ilvLp1t7Oh4yLAjEGufc792ej47U7WQl
YBdFlfUSA0cJlOP9ccXGssgk/0GYRpHgPDF2GU4sDU0tiKaWLqIRp+0WKcinp0f23GxJDxC4BBPk
liz225QoOGEIQEmLfcbvdRMhAV/e26jQRAtRl1Aq5j4ymoWJ8DRAXhvfQFg93JKUdzHb+H5ENr0+
cN3BrYHOFva2rGDsSxEHnVc/udAmCCf0/yio/N7SqvFno0zV178mducaWIz5/uNPrP13H8rB2LY1
vMsGXpAlzBg3I82aaxS5bymSqxgLkjI1DOXoO0KV/IrPB/w22H4ObwDElC28gnCDVZsQ42XiOhDq
BRwoLFD0nSX+CZ8sNVjKUfNkPMmLMimIZ8/L9zVWIjb1whfMD+7rbrR+tQeMuth6fslFmSBGJlLf
KPcjQhXKgBW+mbeshZr1E1vt+H9HQK2VQJbCOv3QhBwBsvkFt5rRFffK2QVpGVNFtFMRRtBddgCy
dOg1hgxjwJXh9Ezj/npO7y+yVQrxurAgyDwUrlHMOs7BEvG+ezXekBN4uH2tVajZ2W2/fTkqfzwJ
7+ISOV1G7McpqVewfDCKTEL6pf2VfthW8Wkha2bi7CSJnTFGFhtH7+Xf3FaY/0GDJ7hcSWMabz3H
bwRuFCOP30i7XOgMqEUBeeJcTMzmXAvbvJ0Nkf7nGo6bKkCWEMOqYO1m2zzlYhUScr+R5BdZ1rom
vgNRxcY5YBiEqhYUMyC4AsuF5N842JMergmfIyJdNAsRphbDv2FAxzZPUCsMouJ3d/TsQl8yCJM7
hwiliRIMI9VxDc6ZJWd5TkFQDtNupQm74VnoJn59Ul9nr5Bd5O3U8froPufikZXI4PR+fUhF7VuV
gApLDGsdS9DqrY/5NPTeuRkUqWTf5BLc7koEwsfhVJ35UN/bHfmvXNRBuV3/ObqGGAF1Wtbs2WBh
faog3iPotDyFJTHngFbHPn7YMx14s+arGqSmsu32OcRAnBv/PW+FPAwM/rfp+7EzTp9EKQJaucP7
bzkVMlnkAl7T4iWmM9zuOGbH3IxTSitfXfyiBAAH5n7k6e2Z9m12iURMkXDTPP/sOUYvOBFNXq+/
0yY/z4iT+CyRhoQCllXmdHDXvHLcD0wN9H3H/gZ6BXFXE11muL0za3xJLZ7IV6HVjqupdJvu4o85
mOj7+H1968Wj3/Nkn7zdWwVXt+K/rNqHuB3HbUsJ5WJjYaDmJo2FFGrtkrUTRMqctRqwp6Qwr5hG
w4RgktCQAe+Z2hN11Ei0+o7EoRWv6Zi4HO99Hohv4sdkRAxq5ZuS/ROiFYb1AqU4EEHlnuY3HiAi
AeLXdJEjl5w8VF8JtyApPyeBkCwQBCI5huqzOujIeDKpZ3ldCvqnZvfufYV9rcvHTYPy/0Tr6bfc
Dz20ot+u4plunUmrNGG5RHcvslGnAcsK5Mc41egAr4JTq7Gcynf+tS0j2NDgFw2jNQxUqfebUttg
an4A2izUwAtdCfPqzyIuAu17eL1EY20FT2e6N+CQTKAbmuhBL31D88USOoX1HxqXFGH74iBJbR0k
3yc7MKM8iG60drE2ecy+A/m5rGTIUkrbY8TQP+KAHkAhn71Zn274O/GtFC6f2C22SshY8Tid7yFW
ccohMY3LwsOqIxT++zhqbug+QaRhji8vDeljI3wg6s545KF0j3agX/UoIA7lxicahD6FSvqet113
DJOeM16ChiJ+f2Q+o6+X/C8eOL0ByUlYZL49K4CFLpymed0EyEV2mYKuMI/zbQtMoJ+mwM2VF3Ql
qYCNqPgM1YxFO29nzr7qTbPFAy4DaaCZ0VKvQqkKqtJsaRAbb6wLusURinCUrKRuv/LxO47zTnzl
UhyE/KhZfdBsrIwM7KdKM+CvRoxXJ0oKepybF23ky8+TMGlXU1J9ETvbcQK8X5syXLkon/MtyQOM
IWxyAkeisQoB/iMqpHsO6G4Ca1w/Z0YBp81MFaOSNPvjUZ7X4rcEji12CYWrTPiCzy6JqqTG7Qfz
NtBpB1rOjh0NU5JffB+dALjHpQTBReJmN+qv6c/1XVjk/NX3vBLRdE4PsfUxBO6TYyvVN/76eBzZ
RxHK4gYIgcPWfoOtlWlD3B9m1xBmklo5SQGp/9QbjxPH7wvIlIeurPT5HIWCTo0K+1HQa73X9Ale
Z5tLZriP+jsMSVuxizimXRAjI79YJnb0KAAP0wjW63BnVEa5E4/Ji/RkQTzdmY5HmxDQtXnPo8lA
Jt3V/x0l0xVCQN3RYWwNd/RtP9HqxP79ClabJnc+M6iFrS9Kj+g0xGIF+iC8v/sTD4cqeej3JHXw
IaA5O7wte8mOPOCHaRiHUirT0TcNqTfAgcRxsRzDkuX9R4+a73muJ8/SzI8SllB64TB4AJbzk6OS
VNRH6Pfb2qlWuM9sPz6CEvkBun1MuBFxx4we3dqyyeJlM6RpAagZF0aSBtmcjfex/37oAz5D9MvU
egXf5UNnIURwSq2lg6RFRkdFl87E8A32sPn4HrSH5wvUZFbk9aBMSJZhMZ/3yzf+7TpFGmgmf6M4
r7x1TG6fFt8V/aGbJ0AjrDC8BJf+NclAvL76klkgy9zaGAVteWsKENmNEBpiSqHe5D4H2Ak3dfSe
Vx74ugU2KHSuoWU9Xl6uYG8gupywP0+ouFttHW31PEsnHz//QpgOxxb/JG7CPzFzoTYIqVYB0dhX
53eBLpX5/m6jai9XzrJ/KY6udzu8rHhPg+6NZNBMLBSOGEcXSsbdfe3apSnEuV1gM+FgDMKKBylo
Ckfdg4j04lEd5F5kVcH6YW+OaQyzbYKUJgvMhKGTEGEZ4rsVdlHXgEt5cdY5AkvH9nkyuOMOt6V+
ZCwI6ui67kpMZ+CLBt7jxGsuvXqdcOU+SjEPK+WvGLW8VyeiAKJC8h5V+9WQ9FFAe676o9SMadei
quwRsyY7uXiW5y+AHb8I9KWma9dddDm51I8YmZFmXNBuxahyA6xTe71BxcPLtn5cKHmfFMscx5CJ
QCO1BhbOlhZCIT82Xh1qjduQG4a6ygfM1Xbx/zPDBmYfWhYQGGlhounWVWVNS2g2hV1a8zK59BAy
OHDE9Rr0kxGT/u6owiarpd4DSA1oq2CTkvSD8z6CVWHaFACuqr5K2uBsd4+p3IFONEIl768Es7/S
aeNodg+fZCqXgM6DJ+298fGWis4bgrLHTS8i9QOl8ww5cPNIPcWhaXjP1PUIdHKGmJY4olp6wbGd
LdnPQsgAztgo86MRrGljbIiV5VCykqec4oxxJsK7D52a/awWxM/05Pziqn9axB8gPZWRBYrKhgJZ
aJzk7Xy6F0i/H06l6i0v2WI9k31fiasOhcf2wn55w9CtM7KtmkXoR+OrxJljefswaGJfIQGSv+Jn
qYpt+r+QMAm6kFogTzUjK7mBq2q62AfA3ga7H4E5FQpCyBCLm8QfuP6Ak90/MFvABXWXqaKo+5lQ
oSdbBnVV8j3Qrouinox6kbTdFpfB1BkoMi4oIGsuzrEuwxCKR8WOswPzyn5Nom8VNyN2Y43Mc8ka
bjSH4JEfQtp9FbuoFMiKaQRwUaO8FH6elwpqgyvJYaWr02BQ8P/53rry5PPWW66C+i650u6pxG+W
HmqbcNHljmeVUKwQFjA8n1VpPjwKgXDuvwynB3gBp/gVmtYK1gwgOVOkS2h4/Ls6V8K7J79GFqqw
2qZdkX5KDJisJTXMUuppW3KmFaY1lP2MPIlqZ4eWvpzURlNCQMkN7xrNR8F8WksEVFzs+B9hm5MJ
8wL/HMvFY7UYz8oKpzmsmvGarv9afDraKRz9ZGoGAFa5xziJJWr7s02wZB47Xd/udr2tDCTe5xa+
B5ItTu8KokdSn3r8ZKqQY2rBZoBDyt0QVsjXv5P49Ko7SYSTjxKqe84k+AmopNo1yfWoHt30aBM6
l8hgINex+bzAuy8Kd/shLRvCKLXydzwUS/RDtjApFgf1Nf3CvJ2rup3ptdOtCLlUMb6xkSHfa/8J
EdiFC0O2tcd70azSigVE7DFjkbONqMAIMeE2P9AfMd2R1nUVbPX/EN1R4+OdCTj6SI9Dc3RXKwnW
LehtCbVhHoBRTkgI07eu6T21PQ/NPvzKIA+PP20aax6GSPDu88q3VaS50ooMGQu/NH1X87FzJmT4
TemI3YzuPRvgb9fo3r7Ejzg1X06krr0L0wgq1Ct5sJsgj3dfJgrTkFMglhYkyLorQyI30tqgS43C
w9OOnuMN7ZcwH884rmnCjBSjpp+OpN6v9Jq1hOagsgRoRnZe90FnE5cJ/pDl3o0K0/SpbL00hPBl
VcJ6ZJ3Jhbidtd71mcksc7Px3yF/veVHxn/wM8j6qZVCZh7j6xWv1f6UE6Tqp/1LYdRkDMaga89G
/5zL3DkgYw9D6I6Sv6dRRhnP6Qzv8y++1+PofFJz425RtihF+vfKYoJuOqZ/o9I6U+Sl5CKUcYLs
eOg4nLZeJPkhY6aEx072RV6m/KzjFf4pHIrNjYwp1qEqMPQFdnpsjKwh6H1pEtuzsI33XvugisBY
Kc53PvU9zyDuPRzmnIiO0lw5tpYQX+QOB22/h9oQRpL5EfkpSggudG/s8clN5dMBbBkGVcFgcEVR
5+52yd3pGbpF/i7iV/3nx8QHAOv+uKLIpuA/xjOcleZ5Elg+S2OTtnRTs5Z9Xd8rGRFIQOqbtjXM
Gs0K0aR16YU2/T/2Wbo6UIxgd5vpX0c1LLqT0fz54isgUvNrAtX5zE9wemUifqm927tUJeVr2AQU
APvHLC+iVsWaQ6bRvv0nCoKrkbS3q3qkjSVY64d+ViVzmeaxQ7ghQ67qCUOSUsa3/7VflLjajqD9
jutob79744vreRs3Uy353GwVBQ1NO8IzpPk0865wk4QdK7wrmToSPWKUmJCqmntFEOACL54PpbEr
/8Bizjui3n19yN0btstMhEESM5BdtoDoM7S0q18xlVKQQpZLY32kCAb6Cjf6bQFitRcKgNVhPFJa
d8LLshV90jwqoM3KjyOLXzus4XuZpthYwWoed4NyXRvHxrEizi57dBEXZNb2xH0C1jsBJJlP+Zkq
fFC7N9fUDTdElldtfBlTwgHZkD0vDf2r93MKPTlAHwFWXqeipp4UCocInHlgbFDH3I65Ppbl+aMD
myJFeuH/YOS3xXVzYlLxxN62BoIzNNwtZYr8MQggWSPgod9cX3wK20O2ax4vPTjdfAaKOSKCX0Wo
kskyTkfuGHOXRIETcf+99wRZPTwgHFiq3SfPrXAztOZN/7pMR2qrG+IWXQNuLK0gejtBZy2vlb6V
nFy0V5aFw35bzqbrVYoG15FniHo9fEoe+t56vI442VKOrNt4mR6Vwu9CdfOwe8vECkcFXPkBTlZ5
mzx4m60B0LBJTe3RMMjtQyPIdH4uJFk1SX0QyXdbqkgWtZ194avqhlqsGqWhShOJfpQVm/xy4ftm
14l8zGqCw3BMjmndADMh4OFLqWV6rNuP3C3qT/epwfVRQG7YK3mNl2mhcNtCuhTpAApfI2VrfEGK
rPd4k7ZIgmdA5k4VL+My4nFySRLKgTe3or9HLYxwqemuaw3C91fZzP5psqC0dWsnSkJ0WHphnMPr
E59J0GFiCovjWO91w+AGgo0W2OE/ElyxZmcn4w71I1elMREqvGGRXesY0XwcRQfOJB3iNDZED++o
dqgGVvuezbqUsYzI3oYhvEKreBKAuh00fjbM2I55SQb76z0PzWkjEtdKCeJJqwTJ+HKYshS0wtii
yWf84MKhcFbKkchMuQJztkm7Lz3H6bzhgFhtuv4TskDEWHL016ASs7J6m7jHL/EHBIueXMb59qu0
6Jwg10XlcLCqwZTwleWvkAJ9+T5Tc7fetdbBcHlcNEx3PnyHAV16SshCnINE+GyFnvXUxHIlKv04
XObHY2SS8xxqOZ3VKWGj1QraIbTPhIIqSTTFotK8bUl/wZgUutU3q0KtHgho2uw4A+xs/KzVcOuX
e3njXuP+rVzzQTAqhY3pSoYoXfJP/kbcCHV40fCNHh80YU+LPNLmw/onPVNF4HuyilA91b3kUBZt
Kbi+EGf3LprxulyUymW3Hq2oWlzYLjCsLZZn2Rqpk02LGcvZrGrVpeSlE3/Y03FVoUpecjzVqEB7
4FtmJJlG51wKTckaxNsyMJkndnJY29K2oYYqib35NQTztzXNceRdhWkTOM6My0qekBX0tgDloVhP
XDIEDhmAXmz0tYaY+AcrPaKxd4wTt0AwR7+5ubI6BLR4+HSmwyYv6p6C0S83JeOhTjk/LA0ieAWX
IO2MH8rSo7CIRF++gcIN9z5QkfcKjTMdSvNUJRLpnFa7ox/i5SV5wQiZP1Lq7WEAnGi96Pji8PI5
co5T5ziJ0bCCHfx/25Z7i3gvW60OLF6+JG2XZKWwg7RU7GEw3sJS2AEUu+lSppB6asxpCmXmJrJ5
aWWubXf6YF+wc5kro2GIrdqc4wRMV6Igh04hTKw07U19l5Y08oy02Q6TEskHGTtc5jKItoVkba9+
+cOwld1K0syL9gIdweCSOvwbUJDgLtIOqFaUBAptUCC5RvRK/YuyL/k9iTcP+wGe0YhY6qUbDX6+
/BqF+VZOFSuZlvqIayPjAoSYhhQ+l6n/cUgS0Jfp+fVM8FU5s+9QCsSq2qVOLm6YyJdXK2PvnhUh
oDiZqAX/q6EX7ctvSTEW86KJRwX4KNzvcpDQZE7lnQ8NRjs5N0XvAhhceEWbkQrUONQGYTWiXqyn
USTTW189KTsJKBSFCAHULvxxBVc47pN9TI0XUXn+5PGWrZ+3O/qw1EZ07HDNWFgkV/kCkV2Xw4Of
Vc/bRJjDeIz/FRO5oB/g5RYydqllkr/aa2+8lMZXJjffrqZO+C3/cuZll65hJOe7rQdQbA6NzEIA
T8q4VVCSoEBg+aBc6OgD38lRx8Etyq0mEn1hy4YmwycPPeXIP3Xs7TftWcN0Hd0ufXqHXwUi3NaE
Xt1SFCbjtB/kiThymPZafPm0IILaKT9/P0n96La4OJ+FTShsXDnyjWp8A1Va0fvE3uLi6vWwAvad
yMNcP+1QaEKCT5GHcupnz58b1ftwu8PvlVWGxx4eIkPHXPoL9hCZRzATico136KrVANTzf8HR/AT
Havu6qZS1oR4FRMSZJwMZhVYsXRmQZ8L8BAu4NZEaLaCrsVJZwhmFV3KY/7E7Y+N73+xZ+oIM0/Z
ibUWXTPxib7cVfQZjPfiD3Sx+qMDqZjPJPqnrQHx6SwDS70d+V//whEt+B27tJUXMw97CxG60sYZ
t1RdH5fUFn8V3/xVxSAWTY8tlFU8q190tN19YxtXoNSkLajGLmqeZtI76DeOE7Fe7IgQq0qpm1Ch
u8lt7DFa88HyWMxeDibjW5NdkcmY+yvc2BhjI1ZErDUif8uOoum6W8GwV9GQNPlLwjEI7zMOL3CQ
8AEUaJCWlPM/+oJrqNyhWguTKwvEXMp380ctisQ7lHuRIefuFoMdPcTycAFmcBpLaXErgMWR4AN2
atT/ZtpQfNCG8bhv4RYCJwg0l8g059MDwjszRiwTy8BFsdTo6fAC72W+GWM5oGDTmyGsn/u1P5vR
6djfSsPzmtHw38r1F2FP5puAJuiqO4wh8GIXOxLDzzQ+7pXf9uH+GW6evvEYaTEdrPyuL3MyW9qp
XFCYHObwjLDOWbXje1Gh25burG6AEXtDSH7WI/DzPEQreU7hknr6UI5XbTXX5qMyidc6YYpHtBFX
+tf9iHL9SYNBwLp4HFe8KM2UUMUFRYKm2ADeyEGH2t8LFyQ6XJ93Jc/mNuvxhkGH5dLzFtx+EnTc
fmnqU9egwCXqmrH5mDUbw8afwJ326G+9uoT5G2kXD1nH80tTdg9dFvip1/43TBAwsy2vTQDDEHr4
mYY6ebN2NbVdSbSk3QNLG3udI1Jff+qnjGKLCCA6HjPjHjMG+XtdGChXXecg+qtfOS2eJ2iTiU+w
yBLWyOpmF55EMNfxpl/BBXt+5LTZUpHZej/aqXdY65fK0AmN+RCzEGlG2A44A9tzJj4JGwuMK52a
WVs5j50/WJrTaLfvyzeVsdG8wfaqIGnX9APrAiGcUpctV1uL+vf94ezR7wOj8KFQbz+8no1Lz/pL
Xn63I9oyj33TIILN+0SrkZlQCnE5eFDq3CmBfOrxeAp+PkA0FZ1BcVL7cyTD+ltOIcNRAi0WjmeD
T4VgW3Xdux2AmgkOuwSJ1a+CcU7iZROSjH/mt9kSm7nep2Nu4eHS4PeyayV8+xzuUvjWTdhm2CXX
jFY69YBoujn4pIyE1pSTx+7DW2n88QUYWsW0yi276ejF8yhTcT5ppNi980yFjMOzT31NQzLoWQxo
peuzWXx3xRGpOtZqsjNkrCxtCHRI+TwEr2gYVMoxTEm2AUxHKKKuxS6Fl37o+JhuOd9HqdT2Q0z2
OTb1FY5w9afTj+yXV//jyY01hJ+1dmBkI+mfVxngj1aPNL65hz2+oWC3BSEvTAqtcqtrm3SiH9OL
G7eGRgBObcHhh7xVzNWI79j5rH9vbvH7H+wRno81dEKAlvOK0/J3cirZvjCuCMblXHCmFd2SCkWr
yx/YT86n8C1NTaOEmlMMqAVxyoxrjS5kL/NOx8UBN72uOD2rr5lSZiSF/Pl5M1/Xz1pbHWxcm0Vb
0XNb6ZYha+2tSlB+jb288hd2uosfoU/9NY4kctqH2MImhMK2ZaNbEqLiwKFOOlz/y5a9GeBAx5OM
jeHyrV+1sVuvdQwjsdE4XRabdGS7KdhPhagHdwbydJP/ptFXzj0Be6C7zRNPPlzMprdTQiBGkJ2E
eYbYpzuG7DqyrkuJq5W6dOPbPidK/NyOFNU3qTbrKvB6ni+eXtPVcYIDcpE2zFDCIVvv69OpwN0P
dT5QIdaYhzM6HG7GN83PsJTafXUz8xksvwyVoQUtV1cnlXepAEvwZE3u0p/EjIP3PqQJnlBUtL5Q
xB8W7t3osg7bjAmzUeL27mUA5h5+k/RCBbBtjBp3jlg30v7wF3dxlWTLXuDWIllVFMrfZJHXWeuW
nPWuzzQvCOplYVemRMNnn6/deWrOdbbZ3gmOwYagZ+fHeWa+N4ZreAZnK2DDui/o2PgnH9QFgfib
16iLHj2dSbNjh20ppvYt43NcdHm6X//VNprDM5jxicROgtjWBk7WwDzWbC52ORvOCar0mg5Atdrp
Jxb2xhG/gRdad7CLC/IyeAel6gMilGDrm0SfgLa/iiuRxV423xKJImpsFPUrZrRScoPORRnykjN7
XRmDb2JvKQFoOqnMrXMErdCcdLZbkiBfzHji9xirYnVavGYio9vITDKMkLhaeBy1lePdiuu+n0dD
Ad5WLLYrGSzVRad0lqQemBKayaVksf3RxyB2BaEbw6s6788v/k4H2c39oAXOcPBmBXrF1O/yFwZj
0BqUDnkGNbX3FLxCSVxrlD7Ak4Yr5WBKRhI9B4iy6pBPeIDFp1VKGa9ujyePOHPnxQ9ltwvxUKfP
j0XlNySXFBmBeeQuLAZTVX3OshBS2k4/GUla773RfFzqbUizX7T6nPTOt+qksAnVqCNicGgs7Dto
FlCdTfmEMdy7EKz17bfTEgTbRQNQ/mTJDZQ/aZih5r5fq65CQw79ZQxTn9H342foUrtO0HMG3pWv
iUQ8Ne7bWdGtaw7GmyCvl3K4fxINOVYwiJA9elE9u4nBskBasPGPoRw/syNfMs667UvBv7bRM0sd
RGUi7ValhmDBPsZrA/yeLEuPgPAOicqrrVY3Syo6UxYW6owKGUyGDLHBz7eO45ltQYzkiM9JmoFk
Wr+JBQQn2SjG2phGtpi4in1+KVHS0ZPNP5i+nGxHeCHsWdJyfPQksQn1eve1v2MIEHgfokzAX6OL
00WII8M2Oh27FgOD81HF0JeJ8jj1NMPNK/D+V/xnakaOBjkP+NmiFa+G1pltM1UbjFOBg5PFUWAy
o+Wu0jiLmne5jO1vtjg8iXBwCDPXIHeze0Ae3i4gqeJi9Td7wJusj451bJDbacD1RYBt9pu72LBJ
uW2YGhiVjFXlXNcE/28BJJhXQaCXhq0hZoPb/bdblL6sKDw1vjsiKoHmtyhSlRAs5jBju6x+itMm
CiSbOIhN9ryJzY2XwiLHVAkQfHqIyeAAXrXik6Mcmppc5bh3auflN9ykxD83aYyMJT5Nx0uWvA4X
NqZgYY5o0qzJfC4JQvsZB3t4lEX12ckCIe3Kcv/SVDS7vhp3YTEWd7HhOGfK0g3kPDCK2cYOV+qf
Am2H+OuxJPSbZNwJl2LFuU/Xakt2MCZ7+uZkNXvRB1emmlOQf60Yhy89UVNPbFcNt0VKtO7VJ8Ya
XrxbQ/9uFZqAvLjoggNodSy4oyvZ8FwZ0UItATHgPB0aE+PE0+kQJU0QtZewTxwihcRcOYv8OLiY
idRET/euF/rofiT7TeZAvjeUXqS+bZc+hObKvDequ1lVAt1zhUFkIC3r/OoV3SaYgCbaM8tD7N09
OGl9bh6p4YikwrF2JPRPdEQ44zLc/k6kGSGQ6mWyx2U8JBXTGrKOoGKnNtANtxrW+G1gUH102Q1Q
NcHORsOAzxTg6NkdKDDZmXVKn9YR/qvWmOPcGQBsDs+IPNoEWgK7Brjjj9OnbQx/Pmnz80zKN3CZ
PxWLxuO72EmvIrB521qXnbPgChKkQ+sc01ANiprFFGK4VIyyV05Im+IEyK2o0rO3gW/8R0fjMBTw
109U+RfVxUYTTq5Pwj7a0urpuPK1Qb+g93x9Hu59rURAx2M0xM+3mHbbUFcV0y93592S7Ab8RWD3
jiSGXBwl1J6RymYnpFOBPZGUatANWsx/18DQMTZbZjjpMOqPe3LxmYf0OJ2YXNIFyVb7ZVeYkq20
5Hz2RngscNUh3HD/LnqGk44VnLLTg6Nj/EfY2W7OzejwvnSt2gbtQWoztRRTnmUn3gtK+czRrFG0
uvyHDWRXr8pWAHu5quboOSIJpgxDTW4DD7j3ztZGwApLhF1PSI2l+DvnQlyhgSau+v04z/Riav7T
bIiMPRtkOcAx63KduKAyUxWjkJubgXwJVfryxevAB4U0zkfqZb0Ry2eIfxstNWQLkuX0gEPCWifW
zoKky8zt0ps1XH7KDiCrhqQ+XY30dnSdn9YbwKI68FlOeRojxY47A9tUx7sGGT2pR+Pgj/wiFUMC
7ioetukTCV+7gquCrLdwUh8Hj87fyxViSc+fbBgL1eCif88nLlVArBQpM/SJtu/ZuCai0bfOGTLz
ax/72wGbVHob5mCKvMjgSadK7XM7UThurt8GjU/49TTrI/S3zDBe8BaQZuW5zulTS+twtZ/soWdR
YoAxWShLJxJuxAsY3KSB0NfbetyDlC3ODKQiPAs9wnuHunOxZOUwXRGFdtUWG5dtnadH62QqRv+I
9IqAZPJJyDnaVba1zTnno95Nn5c8Gr1VrKsuvyUPU+agX8Jm1Qyd2qRLQm53NrhGRKUBR4h7zLec
eDHj39anBFWdr1zJtCjCc70q/oJoijpskYvlWm3j6lexvN960QLhjq8Wg0yNaorbmkuoWrZNt9mO
Sh3eUK9A8jEuRZbEideVWaMSwPycKczOWOSkK7viZdm8BN6xlUjX34c4VcPD1bDxEBlftkxKkqSI
A1s53lZyRS+z+3YQ8jPUlsxw8NzSGv2sHquDua8ODw9SY7Tv42lq0GTuesCxMGV8iJ8hBYiqxgIb
jkbbNDMqfT7X7A4ItasSQUdYVth0ZFcD9bakynGNL+o9WLfbPfy3FSBxmbXgj58J20cKtRtaTdT2
GrcV5JYUmSho6MI4rxkNtzbJLa9z+8NeHLVVQh6KZZOngpRFvGHAWiHdpmLzD6F5od8Ohf3kv1hw
lJEoUMFDYETp0OETAavONfGVy3q6ef3dWOMT/W3ySdH3ENlLR1mZV/I6GKjQVDIUoK6Xb0gwBlBC
fDPolYe0TUO3wLe3LW8N26BpJncx7OTPws102b0Ainj8RMtLOvuBf/xvuj5SFQg85KYhIYk5BnYl
ZBGPbKo8N5ug8B8j95T/qY1HMZl6JjFpmR7nyvAoAENFFwzbSFSS9WneRZRtIxSjT0AVqePhm7yw
j2cMMtjXjmf8z0q7O1rUpYmivracB1T7gKD3y2wwEYuZ0fIXtsuUe+QdXxbmkvRwfKOtxxtlwezR
a37wRYNselPzwoDvMAxHDv+QrKX39StkSs+RHO/V06fIaGkJ+4OtXKc0tiGs3j9atKHRN59ilLE1
xgiRJNLa0QCPoMdje+vA4PmuaWi0tQvXbJLWV4cvCscytjLTDyEHcYnDP57XV3msCq84qhOxyWAS
e6FBhMlURMrU6gnPKDMz/avooPru38tjdiVRzFTq57BAE4T7+tXv0Kq1T1z5vUA212sk+opmnwWq
Gsvp9OQw1GGdDy7UqKS0ZFuYTLNL6/BJ6CgekAy8vcQgE5Kxmkqaq0ZKad5fWRMhLoqP83H8/CVu
ehavgqANF3fPXFBlsL7G8xdWf8B2EkBo55vsQDzs2MO9OHzCqOMEahjrtzaJSwClqk2jZIuu1JL4
X/pA1iQVnHmQlCNzsugknDWi6zwZcgwQF4VJPOWIEDqiY3eJd2vNsDU5qVypFsOZK3ZkfUGsBlap
oX5FSiW6810WA9h9oirR+sDP+kE0WbURRNJRiweYl5SpbCJ7WiHXGBPuxv98jsy3uJ8q+CZoaUge
wQdthwKjSjuBWZdfHKG85IpZ+Iqxim2MSh4iOSYNJnkOEJEiLJ1jghAEOjyDKEnc+yb6rfgCtAIe
PhHmUO0Qe18jQs0jCBXoXVZYlb/oyStnhVYP/BjbzhEqVFRzHAxYRn88ejwI69ZcwezJQfJROIn4
eygFANhBaRx+PigzjPfW/tcIQOnxRnZ6Ns/luDhQxiTgbE7VzGcrwBPepqBwH00Dn8TG4m8eAVLE
bDnJS8xUuokPK8eNAAYJnO/EkbQMAm4P3LsJl78qSPVmsAyfkLpBseONl3t6Hi64CYO460OfLWHA
qs/yg1stsfCSjQpZylsfrlNalhZ3Ta3qnSCCgGhpLzBKXqZf8iN7m3g0KwsrUxB/fGAoc+gw1PCO
/Ddscyv/dTAoumcVfeWefx23M21BSdbRBSz6ELBzgvQiFbQafx9Rzl/SKDrdT/y/D6H+GEWHYqHU
yFaDTHStYdQx5Be3tjtJKvs+iYvHEBuGP2GFCxV6Ha7ifkPu6sKcKGGdmdoO+Be0Kp35e8nnD1VX
OQPfzOpKDutRCKrwkhQzpBzIFXekyU0d7ky3KSVHBIrTfdSeFoAgTzZ9FInqhvMpgfMpFG/cgUzO
DRdYeN/BIFe4zJ9eD0NXdnGXr2t+D25JyIx5nY4L09cqQu3pmLXIb6W5j5/jVm7CYR9efjWLb/i4
ZYBMLHLE6gkhPm/+WmK15BAaqHsn55ETGLUzkWlnBn7K8KdQwRd2Uwh+BQXIVTHviSKrQ1q5O9cd
+q8PA1mdMHKnqUglFph+8A+i50VyxqreAofO3s4Z2T2WdTqzQ5/79OfMKEE483ZL7YM4JTSjrP6x
pdfVdkE7IPJ9FsBQKCdfRrsS8zOWLPBNu5Ep5E/Iw6fpLtfQ9RdLGklKjctV3mkvM2jw5qwqxZRD
CEKqEUO33WuxjLQGFK+BKXPIBLv7IKUsFYOfYHooZn4eDmrmpxQ0yQ1aTH8fQNBdqQH6o5vdgNCY
1cbDMXEiYlwMisapZjiGCKmPmkojyGooYJFVvtOpwa5j7qL3tBXGl4BR8uswrx3sltTEOq7kb8/g
Aq0UXouz2z4tPaMA507ZIvhdxBIeuYOp5f5xbVDjqiQsCePQaiZQCtcQgqT1nUPQid1BCIl2dcTH
sp968x/JMcCcRp3uPYoKwf1Ca6+qZdTHd01mkQmxNwuKG9nl4SDYIohZbN5Y43ufhtwZAKdcmNXu
nTr/BP9b1HmslL4OkIuJtUZ8YIj4OiPbp8g7WnxpIEbP4tBpMNZCgC+pPpINQ1cXHQxhtpFUbQQV
9dadj+69e+NRi8IbNWJOBQsNsJJ3rqMPm+tNYiR5Y9RW7DfGjWTdb8hVRiqyNZO+K1OCCpzbBSs7
1OOF4qzjslFLwt6ZHUNBQqWRW/DK0ilLNHJdJCHaj5V/Zfpub2p7yU7oMEIYZ+vQxz+1nXGF/rpN
RE4nrZUVeSaJtcv0Gx0zv1KjPLGfe5JH425/KrZ/z7IMoQ/fHtzDfvrGnGeifsRtA/7sD1xW/qrD
T9jAsnIGuS2AQ1lDvs8Ru5nNyM6P41Hb/clR3uMx0h9oAiyjbH4QWAarjLYqXJODVNRSCV9aJRar
F2Qdt2ggjxA2gBdhl/aiFwa+MUcC2a0Eji07+0/Q+jXHDUh6CfkQ4y855Hd6RPfBDNMOyQElo83x
VBP/CbqWm39QfxDR6VQW2NflMMOKXAGhgwIQcKazgIBU6S5nnjNwFpG4Ne50h10EAyTA8ksrrd++
3sxlOxa8jgxpu7r/b3KTzfxBtoFvLkOq0xjbnsv2xqCBaDBFb932tsZaJ82nBLF21VF2T7Bw06uw
L1wQLi/6oYsz3bTzljgzf9J/MGeOHy1zhWVAAWETukUSEzNo8Fdzd2nj6pCOqZn2S2abHBdO/nD9
eFim+1N/DLrx/1LN/E5TkJWojDFO2YcQXlltVu3y4yHlubUVTAMtXGfKCjVGaHTt7Lr3nuUu/4LR
uQXgbJ6NzjFIjEkVIFufDxzqDK8aQ9FDzQiKsLrNwmC1fHoNNkosM7ggZ6OVV0wT9QkIllXn7HRC
iQwfP8jOC4c4Buet/Igeg9LPg8pAAk9mltVQQ/g0veXySj9tkk+jQSP33gUl2OudcQpxvlTgIfSR
yTxL23sSV4axDDxfQkeSTFftJIecfp58+lI8HnNteAD+q1MZEWjmWRg8vOt0jLoLUL8o3LGQ7p6A
4Hj/OcoDzB1uCIvLkZ2ZZSb4S/aC6/lr8x5yJ/bz030x7DGL4BAOsRSae4svjaPw4AVTFR0zQlnJ
+6k3d/6eVjDsJen0lEPCL/DrF5uJZXW+BjmaCnU1JMFzQrRA9pPIEDnplbUzD3QZBYXjhlkpH4ZV
qbX3TqsSzXstcxrWUchB3u1f0GjdnhUovpRj+b+WAxdppvRDJP5qNK23clIcOVREzjtFWiRkVGRL
qu0NvRq1L41uDp/3uyo/CMemFSCvSkVQ+B4uqavRcWbBAYr5JOfi9ia0woq4CL5ECSp0rmz6n8RQ
K+mh9fDrBQjkfxuT5XBxiGulGXnIX6/5Nf8Jysb2kb6GV4UFX2bsf/1vbf0q0J2gS2BfPNTdgA7w
fdERnH+GBg0TioSxaCaGBVYLAiAPsLgKkf/5B8Nd8lCZBZvL+97X2ItY6lO3i1DsQXW6qkycTYr0
Ruh2z7464G5TA6NjopRXoiwM5vlQ5iWq4hgkubczx0OKAH4DWAHTx5wdfKgTYbKdHiUiwenftJUG
rt+ri4LhT4xoRWBi8l9jk3w+culr2nmjRuL4euylxIeYyVY3aIGFFEILV8mC6DA1IQe1a4AQhaO3
bXjOkz2eHplNG4MJo8GALPLsp6oJT4lrrh9wn9ngivBTEy6U0gDp6cLTLDWmpAJFo/3GhzLpGnO7
SGFB4Pu9MlhXpsyS9FxbmWxQAjmJX1w/FQ8kOYOsFl8enKywJW7cYbB5j4jxQLC57kOkteiASZl+
YFI7Ti89jMwPInW1R8rXtEk5auWaUjibfYDO4xPeo5o8JrxD2So5Qg2C8liK/baRQ5GBYo2XL8aa
Vkwam5dFZonhsRsXL+QSuww86dc9A1jiMtVGtFw5b3amEja9F/V9sskLiUL0KlXSfwKnX297azBs
2e8zNmJtedl2Msxz3punTEeeqEnbI9u7Vgu2G0Kf3EYRM/F+DNXF6zVAobDhsm6XY7frBT0ZeAue
BNVl21hrqzFb6IJjvrWYGnC9OEwh7RfX8GSQpWlrt+uaT67Oieul8H7qybkA2R3RXpNdWKkgjFjs
kZNRM+NioZDMw0STl4M4NX83ER2fQslLZsL99RJusGuZN5O4DQsiQ15c/UoztbWchLq3cg+kX3ft
Ftxr6YbsEojaYF9+Ddz6JjeCwxooX6c58/q/TnNkbvPGJfPZWowSN9kId56FqpTljAFbZLuVzrAE
CCY1YMNF0U5OXeTKWKbLy8CRaZMdV0pbZ49TPCz8nd8o4nA+sfY/r5hrOwKZ4mRwijYXuGycDtfC
0B+pim9USnVhg4/xCr8vFyUKeB+qOcwCX8vcxYpOEAMzRk7oA6Rpkc2c14f995aiPs5DYQ0DYDks
1AIkX7M37GhrkeoULj07FePAPbczxlEaFESHRmeQitag4jC3HZGkn99UhtF8voi01LbXed4Hxaqs
XXI5eBuMnamRtokDXEUiPyCsEg1wbts45rqb5wRfOtmn5UnIatXKmCMSw4sjDdBGwg/dOGBewTLj
oqzIVXuo0WoVkkvD/T7i+2FHAD4dkwLtlzcAoRSd0Jpp35EZ5K2RzWffmr1fVJ9PMBLM4a7STvzT
X01Cxt6Gm7hg+xG6nN7zsYJgAGlLSOS4NEXg4n5HlfD3n8jpsvohGpOTH3K6o/EU7bw1sSrunVYY
nzmcSzZpC56WsOXfqg2eljz5jbKcDcYFd1JJ+5j73izTDUrRsn5BSt3IYjuXBptWrheuzFvKxaTF
dq1m4eCC5V153kzAc1w8wLWKQ0prdDk7TxMihwaQcaIJzmAgLE1868rl4s+k2iu+IbjXcFwzlMM+
U7VKjmVXvzGQ6s4L/9G4QxUKMGgkZ4QHfmGcmo4pOEy0Oz5SJ5veRyjv8cZWueRZEZ8n8/IMUVv9
e1lQumc/tKWeuxKQMzkCi/Nisc1bS+WM8f2mTyy8Q223+T5OYgFTQq9bsUgvGzDcg0AFM2lLzuVP
wIhA5UnWzVoI5O3QIiFnyVahf1VhHicSpXzB5gMOulVp75LKewofvUO21LQ6bix/neV0X9K1/UAp
lN2d/WX9acYEBa7IaPwlxFlldPPf+dJVoyuANBsQTjFvTaKENMRG/donuKBiydj6Z578ra9J61bq
c3LqwqmbUyI2lvHmswlNbIEyFUjuiM6YwRUjCJPVs7wRUewdwn70ZCqW5whgTthwq7sxjNI/hTos
cwQp6uiXxmbVcDZz3n40UOyRBkv6e+khwSoadP7WUUqntZIag5eQ9AO6z5TxigRTMTpr0xuJM1Iq
S/DIBxI9KTPnuRMlAL3ZGf2I4EvA5+4tGIYCstnskFUeY01Ww7Nv3WpNTlTKfdQhvmaJcfEOk+uW
by0cWg4NuyUaA9P6jCXKWVT+xMVzem5647WAVoSE3fSPnN0JdEGUl1l8WuX9TF9QRYx3q0n5DaYa
eMsg1g9JQM8GrPCNCnC+KqCZK8vwv6utKnI06/n1rkDsAcN9UQdgaBWDi70FMiOayZZ9yxRv8Rtd
DAAQUmihdPRxoqUxtqDitkPZ2R4OYCsew+Sxs2smj0e+JHKbj1NRVtdB/ZZQSHTB9XH1TmHN5g+s
WuDzygldIjuoruGnMcaV1R7REeG8Z5zPbhNtFdeuwCff4g97IPy0au/LdJm7VwH+Hw2A6vspklfZ
6Yp9tdoFwup8JLJwmTk7Rch2WVhpuxHPfg9Nrm0t282a1ay3vdsAgOfSbYGW5MLUKzoO+O4/OU+A
4MeaBKCtef3Y8/RZNkUtfz77vqJoCPWCTu8ReD51gPQrRrk6m8PDuKHdoBY5hMUhiVN8coLKGHfg
+IMWcEdA9tLBEn8HTmIne6kvelpQQm+K8b/KITHzPxv4OCXOE7TWJo0YpVxpj81Hi9kKPJYXi1Qe
ZWCnLU1683gFL1Rq+XGqcpkfx9TBFwOTyQ9xi85vlJO/KZIo/k5ZpJ+yolNGUiJsqX0GMABFtd7a
HyiheEGxQE0ctxzCJuVJKEmqT9250cTQ+TcfwJsZqlLCsQaXYowHEYS/TuIYjApqF07TQqPSg5um
QwmJfF81Srmbpl7LABvw6webXxr2J9sMtrO8K6nVo3gQ8PGIRoPpaIz9zcvqn25+cY0PQYtI11Dv
i0S4xANjGXm3ms1jdM1dKzx/nPn3TxPE1S2bznIo7WpcjjXkqys1ff4DOPUOTLD6unsgtIg1jAMg
qy0OsjbDf/VYPb6ksBnIfYPFWH+xF0RN0a39hyz5g7b5MHtQzUiXCrvl76x//RoikjqbRaEJY9OV
0sZ580VUpmVqs/IvA1x25G5qlwrWrWJL9ETrtXegQRynlbBqosu4mfCZGVQysP+0T6lk96pJcbPX
8dEuIUSrh6/gICbTfeY6U4ZW2Fu6YXDpulHSvzN8Yx3vIHhgiSi8rbp1nk6rxnoyK8bpg1nLl9eS
EhAJJIm60cPn5o/wchm2HyMm8YNjlpMRBYF74sUFfF6Be6tChGvPzuFNbkVXOov1PIjWvEh3qPnp
F/JUl88sZjaNP1gUcDZKGRklAbtOFQXXbQhMPk6aHYE9CuCqz9n9ihNkDJRLIvDwrJ8kwV6SvOAm
pdU/gMLq4bSZ4U/wbo5igdfKvy/WCjV8sTghBUvyHaN3+x39VOEdx994wg7O+PBqbaIbsQ30TA7n
pB6iQcoRlecaO1AggtN6U+2Y3HqCrl2QBbnD1nVkZrkQv/VybU45wlWQpLgdNiq0F4+Yt385nf20
w2iADmUkjY3FyHDmpsNPWPmEIpFCfmhjFEQTvNSd7FEG7rNO7wXVXLNNel1a82anL9LHA8GMjby4
D6snTA8Pq4s/Kktt0aFq12oAuvAeSnmC1lMVqpnxyhVSBLX74ux5xHQA9jvCHLYkNZdmrzHWrDa1
DACgjQXe9fIjYfaXU2ICOuPcxqUF47TWx5lPXMM6HixXWcye01ACr68joWL7Px5BLyFI9kzz8dWR
M4YqCtjZe018/mQpNYdZIRQQ7/EY4/kS+/CoOz+mmoO7DKjiFzo7P0PTV/UyMVunpCdco6WF/Xng
cIM69oCxoOriOd6GwLGOY7G5hEajDQnI+J1O2ykP7lxxNfu3s1Pe6+riYPQz7m6KkZSLrUtfWKmk
5KOlxvxsHudG0yr5w85gf0skGLlMwqjAEEbqjnfqG4EAFW86UguzvxJ4vZ/kqn2aIWw7SlKSc49b
dLeICokMY94BOFc410ZH8rud6aSyMsBC58xLeUw0M3qrmLca+hWRoIOTSA/clpfntS+YdbgyFDRP
+87bIGJDw4FAkmz4wEPmeGWYThp2zU+GnmKQg3rmK8T4OlnGVlkcIqxYOKhUP0gOE5FLj4zYzjEm
kOx2tCRFMaKbQKmg84qRm0e0pR2UmxTee5A04KmonMA3i99bTR5dARSdM3PReMbXUMB4secsuBOZ
nKrcdExEbsmuXxf7x3HBe4aQ11jsbKqLG99Qs17BbYCTqMG1IN6Bu72Q8fpYMyu1NIry8qHaP1cw
92FX5NVNzi+uCy1SZScYV1+sDgRr6EkNWnf3V48IPUC0PJwiA4dhLFrZG37MYz/4E+p4b53Jw/oN
SkDNyitdk64kohrht9F875bqymX174/gWvnt4gXwHf/1zBWt35f1BNDcZdKis4tss7PvaPqEgNwr
NHvLKAiYBRfCRZ+ttNM8sWMLYg4feQd0za9XoErITDj5AQYaJUrRlWk04JwqJcq7HU/vLRZlNWj5
ecRn5h5N379NclXD27hFOq2cidURM6NWnLM353l+o3Eje5eVx0RHvABVO68d/e6tyw89jlJ5MiFL
3sR1vKxK7jMCgUK4W+V+w1Tm/s57iztaqWVys8lc9qTuOHrGcGcObHasRJ4lAyhAILMNr37XomP/
ItP5qDiAe+L9H92jDIC1ZyqfJ8FAiBxB6skxHp1hgycxKGRW4ikbdth+OG4yjNKp9DH0dx+jJzmn
QVAlH6MRQR/VJNhFznEQNlAV+Sdg+zKCzrW/52LRFzpHRnuS7b3hise/rN16kpPyaEkuj2GMEdPR
RXuZZ/q5FhiE+lr5gm/69fKmvI5/c1bz5nfqu9p4N69NqPWqNqZOfrFLgR3mzUZwU3Zr+ZIQ60Z7
9NUpPkac910m0jA0I6p9ogtsXat+HGNJX8+TyR7+TxdagNoN0lV8F76dawfa6hd9J9r02Q4nfm26
1Z76N5iDzI0Wz7liLYFztXzCP05sCXiuczxmYK7hUCJ9FFzLc/z1Zt/sL8co3yj+Ekvkrj6JmXSJ
FkKmy/L1JqTR+6LD0DpX2pGSKo0q+/cL3fRGzE+oUnxUIjh0mwYILxhQr2lC2BxDiY1iyubC4DP3
G/CAvO82DLn9Q3mwiW2ooioq0G91FN1is5tbmX5EJ9V3rNf7TOq1AwWANUhbH48bBM82bRKMN2+0
i/aV5CHpzbzGJyfn0zg6toC2lmsW2aTBP+8IYKi/HlDCwQAwqOIaCiGnvfomb6x00/9geB1fFzU7
/oepiQp53Kp3wQ99CjQzZ7lPrV/MVbf2TNxa2FLGIphX95TjjFK46jOQr9MZS/iFnlVPji6oo4Ti
180wFTKIy3OSIahcC4JNJyP+g+h84RAwAAAR8AZxJskmZiUrB2ad9wqmeyScx2SUaLOuKEB5cnOj
N3kWLwXQWmBoUSlf8CcpYRbPaNfwicTXaClT34l1fJZNR9N3ka2Hd90v2UwAdZWkRJdmRj1S2Aln
xP8ex+J0+f4mDhthkzTHsM820FM2ZH6G8+nvVr/bGqi7YN1DemSENUwvnZSZ0RXcEMYGhU39gHyM
7+YZG6WTO4WIVyKaxD8sZ5TKkUN+uvf2gFCFch+vaAyXHoIKqouXY54KLGC3872u8bzENPVAYHat
WYOb7RM37z80ZHPM4Gaj8SykY2SFGbwKIWBc2nwLEOIZUP496Gdcz6PEgjzX+INKgI2gPmWhCI05
vj2DXE4Rd96rgURm6CJihFmoPGFJSOrKX2PbTHEs6gk7oVMznMCi0lcVrbEGQtyi4/o9A0vEmtiY
fXm4wbpbY9jToGhlB5JE7b8gsaXSw+S4+5TjTPgQYehgWlexwTMsvJ5uBd+F8GRN39LnpvC1pKOi
Ngm2M4YMH4nfLe3b9nuHuGHsrnTSbj37uTm+pv0FhB1l6Jc4Y2SaYU7nxlWGgi2vag+zob5L3BZd
Xxm5bJrxMYhnY63nXh3U1/rZuw/5wPsEzB1GZ1X6cIW4640q0cnute4dCHpyRa+EJ/g0v6lZ+Us4
adM+XtMJqfgHZ2CwnXvtKnZKkjrFRVgBQydfL0NniUpnClomLzT2HwG8FdJMfwPUSH6VHBSOK5ff
vhYAdnjWthzUFI7Xzq0Y7WgA9TTDUeHy1Cbv4QBUwe4XGonnGHlzwcvhZt7En/UejKiD4Qw3AyXW
qw82sDL6uJIK1b2nTrQS7ENxLZ7y0C8CM37Sf/5m6d8QshAKZcLIvKfcAU9DNzXtbgwmLgsDmexD
xgjepUFTEQt67aqCaMJQSgpfn29/BJgrdYeKoGjobvKAcQgrcyQchOCo0el8d1nfsh7zsOCOEvr+
szmRD9q4AHrq19JouUh45Y3T2vQkzCRRyl0QSEUOCGXvm2CNfCw+reTEoDe4twUwpaZPt0bxkOaN
6RNJLR7GPLzBCeS9ek7+05SMxq7TYOIQC0Z2FhburV8+7ovSZ7VcRRIBjP3db7YNP9Eyec5eJaZ0
SFIviCq+N4T4cpxsoU56VyJI1B9lV98NbVqPqye15OC+hsgCKoj0BS68UsA1bwKzM5HKU7KEn8Cz
rnPoJwo2Au+Qom6nWNQpgVl29COOxtlXr3uuBoN4UKU63NJEe6uY9+Qvcln01CThGMl1lJ0+Ut7i
27ukSVGHuswFGiaqxU4JA56dUPV1/nZKSr+c8mkFQKVcZWcCmHXTUXtflRLOq5HcZOP8JZCUMsYe
2gDY3uDsdWC1NRYBxiPW3I0lJ0J3kmRD/hzxyjXevnaOZnsIqT2D6THqIHmEntUuStYwiuUuni4j
wIBwGQFAcyEpKWfe1bYMO/mThDAEQWE6WVKd9l7dfKFODM9raRAg7I4nM1RhSCmM4jMRQSaIsrz/
UUttelOomX5PEbOaMnbIMsrNiTmU/lzGEuOduYD1AJscJUAXdJOBlAWNB6N/aWKju0+5AlEnuk/A
ZM+4bj6YQI11KMr42lJM25xK3I7nH5RQpY5fVaSclyv9b3oP/9aNxoC52NjPEZCNhtkuRVtAa5El
m3HcC73E4pvMiHu7WMoJj+0a9X99pKUnG3ui0YO74+xnf6dm3lK7mgzGcrJbwal5qwz24YBsGlZd
F/l1Es4iQ/03NtioISoQlQHFIM7nVV44TH+PD6hyGVC8DpuWOiQ0U0ZRvr1JNkfqM0b9Q68wNCZi
1wEw8Hwc9iggYioiK7emIyHxvJq/pFu9CCzWb+B6ZdqRk3kAkCO0o32RVOk3HvCLvM5sJXr4fHME
JZ0OhYoQ3V3VRhrnU0pkHh1LUtZEShyCD8glOfvjbdY+jPVwjqlsXnOIYa2D2biFQxHl1pC6U66J
N12AfMbvRqKx+qQFU5yTOetZPLv7KU/4sZIAGoOspO6GD0JlJob/hQyF7JETb0Af69FFWfP1GAnr
P20H8crnxZcACrY8oNaRK5fj8l52zkjj0X0tRZ7cVxgCnxclQxdSHIjhZAWKajNV7D7SxKmkiPjC
z1HKK5TldclF9975z34IWqakNFJD3hEHkEvK3PZhIEKTwHX8C1W+fCeCpEryB6eQKYoPUCizgump
gmmk6JcWnU+nONXStVWQqyGz4CjFLxOa9nyAexvDXDnJJKlqVkXvTAZdfupxKOEA6HDn7Fy7spD8
6AWdABd5u/b/t6D8Z9rAPgKK2cWMUZ4htsCuiwXdg0k6mDAfiasU1oH6tx4Nj1kTzqmxRTVrVqxj
x5sn1QrC+5uf93agwzeecwq6vVFUVvHDQeWcOmqqteK62lkl9tH1UpiBriIifK6AFYY3fjxdX/is
0fcGNs42Yuh9Ka1gylp1n9Z7mRBSsYTWpghpO9KMkqzjeqxdXmVdre0YMFa8lTziMUxTVdFU0HJI
yV9ZSBuHhzcmhsP2Euqt4Z3zi3ijYFv1+a1oxMBIfVRql6hmQ3h3MwrxzwYSrXmbUlPeEsD/AhGC
aHZDu3yc1T/ZcksgSzOD72dMspEXglnygqzQrY0v74O53INC7KahfqVc36OurMVKEh1rNWEC4ZGS
66JtLKzGE9ZmVqtuf9qWvJjbLrcHri+w91ca4dv2q3O40d5FlacOxS91/8p9cgz1VGkrz1EyCsA9
HY4zNvqHX6kNmKCSA5iSlsgDJEV/uT5TAkUfNAg5ilty7kxTBxQMKz1VmUmS96/yQ0xYKKE20Er9
TjODe19Nk4ggpNjC99Qn+XmgoXtpBIxIRCuuMsdJo/9w9Jo2g5RmPIMZHVIq+2cFdMO79TSL6PoH
fjAjjKvd3DRaR5p/sfpFfUYuZofQWTLDxgIlHQyRMteH0JQFeIEFE1MjvfyQd9Zxb8xBmWr+D4Kd
7JFJBIJvp6qEOf8jkz1hqhoYixpBPzYBpOdAeOZJEPqc3Ahs11FQpA543RU4Owyfy1TuFrVV2vmb
ao0BabDFBX375SJJmIP4Fp3iQ1gt86/QndjDlI/ThZZPJBcFlxpv7YEdXkbQk29Roaa6TzXO2jEt
T7ttDYIqWSrB32m6VwvdEOP9sR8lCRRuDZnbeAey4wIPbhqOxSrXc7fjNmX3AmM1YHvs92CBXImA
jkLIL21EWNUibkAtZV7G8QCVZyIjOAfI95MdtISUeDjG90diejoS3SGamgDFTNBuMeONlVn17km7
Av8ssVykhwNSQBVEMOiLpxd9o7FBNyve4ktkrZ1ZtokcFVL4vsyWM3M2gY8optBgCEcOnLO6CqIO
n7saZX7sIm4NUtDpz8gOFQ6EKKa4OBW+sJZ1pNj6SexhKef9jQoj6L+lxZVSXp9FBCFkBvH6xLhh
X0n+t/LQEaUjSm70SaP2N+s8IgNFQ/e0RLQxuSwkTk+ySnNEXM1I9ZNMI+3wuedHLmkoq0QWuE15
9lezFby95mjp0QJ3u2Ap7XVdbipqMfarDHFIx2Foa9KsO4CkaETt9Z5JaW0kcBj276nTi/biO17J
U83MKC+cVQNpJ/kNJHxFxfg2oa2DYLdGbuuM5oKbEyccjUuAMwjJ9MkdsP6OADiNuiEE5YSvhxOj
ccJCTuVMg9NLDdUa3mmycUYGby+Gl0fIkgY1brMCwREqxjOe+JMcRsq1LJOxRglMnNn+/GCBXQsY
XsLeq/ohsJmwnhULUzNfhufNdFXMk81ed8FcCicCyOtwaQPVhuXnUb2raCs0/E+3DUr9xGkFxXBo
QqeiWbFj2enZZ5CtzdOp+jXkTsjIjMVIq8uoZChd7dL4j1cJzw17cOMQurx300wwR6MkLYplF8++
tcThu5vvWxhoy9Dx87GWXBnyucNjd6tlPRhLqD/yVCLPm7JTuxwnCnW/wtydZpL8LnGNm3Mgw0vR
qK92GNqiGY9mVS9aY6og68LK9oTbKLHV7w760DMqf8y5kihNm1tW00fG3TXMdMFncYRIE66T2aV1
mq9UeXEODd+TPBJ+fLPGXqtFvBHFZ9IqDIvAak15UBjjjH9FjNV31XYfRGt9agGzkOeDz/8lQ8fQ
Gf1+Bf8dnJMMkfjueWkg/RAMSk7yBfqMn2L7YNDbNDmoBE9qNbH9/kitR4y05naXNBJebGyuLMH3
9gVpwM7ZFxMs+kgEO4GHSWnBKgGV+YErx2ROck5Q/RCvSoLWopgX8cE8/EAPxhM8LH0reGeovYJS
nkWXac3M5s+NYnAzaXyQPV1jKZO/6QfyUuzDxAw47zk1MPDtNzgVS1JOAV9xkAJxINBhCrqlsDFv
+e5YMgc/ljVV6pOn9/qPQggnVYE8SVJLptkCAz0ZvjtSIlQRO5hMDdFrNnH9Wla7kDp1I2+CeGqq
Maaqt5KhqPFxdUF3bmJSkUrEzZ4QQFnvkFj2dTPc0uuLItx8UfBAeeuy9khO3MCbvMGfes1pVExY
KdFmsua0uz6GuazsxzUQxOuoEeO1Avi8qrU6JsLwZMGu3zSpx9LkfTxCczdN4CcbfjEFzm7ySfxM
7IxBWdXNxJZkHaG4o3KVxpvUcCk88tkS13V1+HZzEr1tHydcqZvv7YX/8VKHvSe3C3IXcv1N1Phh
U1aO1vlUrbgPOjCF+5h4duIQophVWvAA/Hz7RppG7x1Ku8EJGnY/vPOEtfPBlWJJ09BiZRjT5UF1
Wftw9DOR8R3zPStW08DxAryNkBNLmA+Rip/gJMVWfBPFH+VxuyrW+fo/IBGnvT0IT8EoLGSlKxWR
0bK1oWGDDcRsocJgxNUF/zF0C9TebIV2vaQ4FFfDFZK3Y/Mf1+TKGEp/rLgQ3ov4NHSUx4p9CjFa
9AbSE4q3/KzEh9NWnxK/wAPCkJJ0e1vN4Uk/qmUrLNDxu5BjnDBF/CMpPOcX36BdvVTy/lay03IN
Y01tMwKoE1bNzTM9UGlQRXaKyZ4OrIOYsEd6DG3aWQkmZ5bJCFTMRz9ans/XeRcyrb1BwToIgK0K
ON2dm895ed1utMZpmc9X+tigqSHdmkyo3JFkl5nJhANu1J5l6dW/1p3zSCocR8chopp+V2nbUbBz
qqxASUSk5d4fR9gTkhJaelvE3JYE83SyvINbSdaB9THJloJGs8hxxb0p4tQJ9GKZFSaHgf//EizV
QRVHFp/8rTlxcBY3vmXB49akOcXwPfbbIMz4WYpNHauByGdC+2Fuo15dQ4BHHpKrSaNZk4ADKDWy
1EkBxB//zV0PYhZLzJHRUWSH7909HvpaehQJ0rTPWzdO3oD8A7vjGKNmPAQZLHtiZjLPX34vdtyt
J5+yZlz4NyEry/jJIuWc5bQkP4uUQr6PlLgc7wvRY1YmxMLWtt/79A8byLAJoNVtHWBIDo1mtmoL
7dH00Z9Ap6zgtcsiY2aLU+FBS+jYUavAu2MJfkJJ+cRjHP5SY36AdnUOoeJRiU+kyjC7PBcSCjMi
hyHxUMfxUHXIzHXqwvgzElj9/pvVPLsgdCLrUE/h2p+KSnqpMufqlFNJJxkp6RMtpTGAE/Yqiw5O
VkNSEU5htbqM/ex+qoINIMYA7RNsFQDdJDH3yQE/eD8/LuoDI8zaGnp1DkS9XuJ+5QRu85FB9jF5
WZAKJaUKaCOPtExG3j984jIAbf9mGC3udtMG1rcV/bHac8i9wRQe+MBYJa+BjI5WXvhkP3vuEsRv
xSo0CIy+Q18KBSvPC135A3fRGd9ZIeFLU395sAO76wPLQTxxv7bzS8I2zkxrqZEoMEQfztW3eSpJ
Fr/z16VzfrnEMNhw2SOGtsBC3cjb8UWNBK19LSiHfc8cYmqWhp7pktkAYfaCG+5N6gFzH0c/9YsP
bUKZ8iq5ZTzg0zhajiTO+bbD50lHDignFoXhrA+Y2DJ5/48DIp4l5qmteNgNwlywLkodsz6VPnnr
XpjXZlzVMfkGDgI4Ke8+BBem14vtjgw1BZ84/NiDD3yYRynHHK5R4DMblm/K2OPcl9FU9RDDENRH
ANJH6gXvluCIMw4HsunbiJoLEtbhD1KXrdRQGEqHYCjmZCPOEkMFvdcc8Odul406neg39vEwd3p4
j6QLitQDtWBWP13RuY7cdk0Ax5pf8vUA/iaZGjIWR3vaHMUKJnZVz/KLw+QetaSCzcrLo8ICy5BI
AjKafrfm3NmKrN2vR9DQoYJdX3L+Qo8Ue8oH70eTIELHJJOe1V4DKELrfDIWBgTolBg4EGk446Eg
FnSxHOQQyHScD2G8na6k4I4QTjoCQGwNCCUzJamXRXudyCpvhReOpZzVlylqsWu8o3A13d0rRm0U
ak9VrqMm8iPSWWJ7XgE76UfyNoL95gMK+c4Mli0To4SSEg47/JfMA2EW5lDer+tiygtNgm68MKFy
Qt2XCXjvY0lV3EhtDrUzSZ1lzH7jezNtVl6Rj/OEfsBpLTcjQ9C5XRk4q9QA8VuLf5i2+IebxdHY
0XdW+brUlpY+c2F4AVr46Lad+MDgbPQZ0cLlBIya4rFghbdKz9E0hPZL4dIz4N97ylqe1kfis0YU
XETORI8EO3GdHMo8c+d/nHl4JS1wGc/kggH8c3tsxik67gfLYbUEp2qPF2SnpS0tVoncmUCwgJx6
vOcYlNMMGIcm/e3/rW+U85uC8tpKj7eUHU5bT6YXpfg8g+5bupFSOGzbkMmwPVDGmzg+6oFvc8Dh
j/hZju/bp0g6ThcHJUt/doEy/5cyC1bMrCcl8trwJES8SzO6/sZn/7sKTw+4Lz+Q3ltOTMLCAF/Q
/i398x+rhjhvOr5fmNcwzU7bp0HLXVWmBZinENIbB7EgL94OButk4U8Mm4VwBqFmizPJlctc5TTc
I1QeoHfv3SBG+rK04hCdj99mQfGWikDlR2dzeh5cpIPPpAiHpJIOwRTza/EPSrcNDEZtK6q0EWg2
0TNEZW5nAWwRjAchcklOVDBbf0q3sHJMJtoewGtE/LvCzEV9ioYB3WP4YfGgbC3bpQzVcA09ZFmE
0qfjBpf3qvWQ378TpavRulEJpNgo6uP0galZgkT9dBBZhx+9JHVjfIW3OCUj1RsG8/fYzhOp7UdG
72im/urqt3z3hdzlefHMbSbq0gXXUGysg+vRQTwNE2vyiXnjX8PjH5oznZEVEocyIkCM+x7MOzFv
EeQ3Xm6XirhBpRRdmgJRb7xxmi1KxiRXox+gSNMeog9vFuy3wnJ99AcyYlglrn+hHSv5aCHGAvGw
/MvxFo/QJsAdJEhqJZkZgbuajmgZezRWc60ICy+Xk27CkjaYBCM4jPxzYPaNHFcf2XgPDLzS3mYV
lrkky5RkutCT24EkBTDciHlIuySFPaa8wuGAOKI+hkdPorRPbReuWKlJSy5FPKvdnRW2NjnMEDnv
Yl/rWVyz2jtK4SSEw9SECAcU5wTG3X2J7KQyjKEW4axtMm/R/1pnI55NibCP55E0yyfgSnUOcD9s
xJrBeQVV+c4Ch7YzIR7+MCkJb8HLuq/DpmUNmbv0SrniROlSO7C8qhZfFkA6s86HMupLxsLEk45Y
XefTLTon1PZxLnCCbgT8nbcBOkKp7xHUI71FEJNEFxENvdyHyCtXwjMqhCpCbSn1815pbbTcIu8f
qgbdzfWzxI0W2XCOgP0uOD+YLKaLz++PRiJ9ClYGBxnmYOGgNdC8d/FM9eqJlLxqkO3HE0dMPw0L
oS9uYvAnBWxKzB+6pmtDdGENyWGGqRDSYGrdC2ImREUxHDQrozQJkYVcd3n+5vtT/M66fPLuFFNp
7ZiXKOVYgE+OLdL0iRX3Cf1vdi6FNh1+KoC7a9xYDta4ZDOZw0kp2+xvhDgMtkPFrpOl4FRNY/io
h61QXc4FS7V8H0FUH3cpDhv69Oc4QiKBk+soiKAIxhUK3dJQ4oC/SJlxJB1JV4Fhmo4uOly2hWjj
gYfGob/F2XZBEMobQ+mTJTKEtSGqjEuc4dKDXsakxGYRlY8NuUgg0vwRO8qhgpsu6kTHSl4bhaez
24CTtAFyQCLmgzyEoRq48l0EQvJcwcaqWraeXW53MBk+eZvKHZ1/v8p9A4thZLcV/AaYB4entYV2
DPocJEOF0tSFfsVHDN20fMysld/r+iO2KJOi8txG78BJNkT0AEz7DU0ergyywagl9QbhLyLfdIcc
+0QEovoKrNLJrHjc8zRHb6pUHcS0CGAJf/1ki9Ke7Y5C3B+t0nOfU+j1v7/iOAjtxd40WN4PJwNw
sa8ekxvuunruDDQWlsAgaPKt63zpu7/1kgwUtpuYIqm9Fhdi990mlk6MNHRZ/u3Cc0TbC7TDQ5HQ
vSqawRuA/wT30ktBXXDOe23pjc9Kq1t9+rkXH+5C2KFXY5tiFyZS8sEn2M5sk9v4UkgSUaM0M9n6
xr/fHRj/x/ebOmMpGQySn/aWhbDU9R5jRIAkjIOWnXa1YfPeFpGF+prAoKFo2cTaxDqRhvlGsvtS
QM29var3727zar5bjp/8ghg+mlqdjNiwC0rvEmjXi9ZSkXT3toZGyRtZGDoDFPhsut4nMPQCZZKS
nTINdFIApZVozB7+JKV6/qDXX5QIzLhm3XHRMaDRQYXTo7aoDwLcAHtN9nFVty1rPpMlTRtHJJhd
CJJgOwCJqH1DMcC5xa8DJrx7ZNQ1gGROovvD4QWtZ2V7V1Hm/tA5lgwTRfQZSnJc0wU1iW01tksQ
RlJGo2jxOCdN8d/EQjh3dryRLuHWnU5ClRbYFyV/DXsM5wWh7S6RcFM7ojsMfEmGdjt1p5MJuW5b
J0PrKVoaL2fmksHauxg+v5yTHDoLh/G2FnuDF8jVhkDUFUFpCRnv21hYAEsPrODduBwmt18L9T/g
vq/tYjpuvBEK4DiTr57y63HYC+g0TAccX2T97KqnU+EUG3ICil5d8w+GqcBUj/PONyrwIKVzjoYm
JsThEk7g4SE7V5rHezaAPYfWErNBP/hxsQfYxL7mUzE32Xa4BGuCgWX/NlhsliyYqL9A43Ngw/J5
uBPsNMdZDVw2oPXDnIx15TZEahZFs/Qy2QoFGXkOUe4AuqEQPF/MfCwmwqBDQvi1bvPYttwXxAp7
WvIJajOwEm+tp9SM0OwdSkJOwB9F3UVrqxbNWWO6tBw3HBntbWr7QLmaE/Mb0KC5ZTUC7R9yP1EU
CDiK51A6Oy/q9GPc30FZoutWv9XxAP9DeOJj314BUA3USaG5lZKqa4UPGa3fcW6GvBp4XnzJbfMh
FJYN54V7O33XwCQc5NmjpTWNEgbEc33CBwFNXFF+aTqkoKNdT1qASD/a1mMBIxOARv0QcsacLt5d
fGP8+TPIXAZ+FAFRHpbFZS1zdBq59/HtD71U6O2rN+CqVr8ExInBljv32zjdstfTniAdFhDFa7QM
q8qo61uMPdSWSMJhE5QUmHSzFDUaOqy7OzN9kpj08Hx/t4jIljK2xShSLAsP1VHzMw1HeqzL3okI
jeXJoTu7JUJAiq9cnwCqQkgE4CcrYhhk+fsKsgGQO7MmcJlQlj6bXF0RfhbcpomkUf4WjHor9iUv
eWZ7patdAz+jZQTkYfEQlTapnaktLffGKq1R1X3sYxWB68EtZhGAr9W+5zvpsDQLo3S1TwWBoEbQ
+ZixQZAXPpXLQuX2B7/JMwvuYN6fgBtkfLn/uncUjc4OweCXVHOD8YU0DwjPULldiDCcSX1MsPGX
rQdWFMG57LL3h3nv+s+hqQFq+1G3rlNdMlqSizuXVoe7sWLlDBi2b8aA8J2Jy0TRxBNdhzViLreA
mZAhRbo81j6J06QVpEloLIMQk4pxS/ijTuh0ao9iqbukZxnhO+IW6VP1L3cujuhF/hiOX/Yhkmn9
GgPV/kZOjZHQRu5gMGf3wl4VBF5EQeIaLIjaYmolqgbyYdNkszPP9lFqH8LuccKKGDaEFrnQ0WRu
tF402m7dEdhy1NItxO7EYDV33fjsiQh6Pe08LkzisGO3TVz4g70kJb3Tl2w8I7c/kuoBUNhX52ve
jQshOIbbrdsnfU/5V4VyzQGoIaWxGmgeN//8X5s2Oszwv2NebwXAly0LrgL39Fqtpg/pcEQH+Nh7
Ar4DPeoiKU/FbD+D6KvSJUYKvwqV7yqN2PeOWKJ5DwKIwfJ1XyzNDLJg2rFCFDn5Oxd3pvJQSU2v
hVPiWj8YyLxJLxSA2TNALHh3ImtuKNYzL98Cj84vskZiK2DteQYgbKAwxvDbItSAKGpDHbxCo4Qv
kWssue13w0LnQbfOJHNYzxmKu0Z1y5QT5LTlay98c/x3uA5yRc7Ze5B+qF6uqHuG7Vx9UmixVe1R
rY4wc2XUEtsC+atnPhURdYYLX4uPv+Ky1Z1WMSEBP4KsCMJcFJWngGLVMD3LnXD1Mb8cMwmGN0Jn
8WXUHg4NA6ezJNe9qNTITHDyJ+aGJ32XmZz1ZGCWYD73dAIXUq+MFzeWj8OQzReWcJZLT4PV4rb9
pfmKpllOkF/cKRIVBZb+w6JFdM/19RKK74QI0M58bCbwF12OAWclHjDBbj+rhQ8J1BgZk4dxNvkX
e25ogOc0J9t6xc8s5wNRvcMQ9+hViK50LOervBLJWhE1g7B+1gPuICTgzijhPZqFTfj4cXPYNvKq
xn/vDx7aLAZJaZpyudsdSQzYtAXx5IF8jMUxMZozZ3sbJWkn0+QIzw/rvcG2PDRovvwm+KF9LCS7
NYScJ/oK73N2TrLSfjysEkVw0q1PTa0hJabQZX4+S681bK00qOgffFnAFb6aVL+3fU74bUqUbz0D
CWHWsidwvAEQtAsZS9iQg0/cl4UEix1tUXdZQ5oTrQm3gd0YMPZEhwaOjRIyT1OAnv3GnWEgsWqI
V2FNimrOyO2CSIaMDABkfaTru1Xu9BIt2I63ER+ZaXCnRNtQjDELtpf2KkM0eRWuNGte8b+xMCTS
e7Qo2mOxVI6YjJMhp8N3wy2eWA/VGPeW2KSJlJsC6L553PSJf/qBIbfVVN4mqPklhU4nUrY/kRso
dPVqLvjVC4R3OuaMlfh3HUFFB1mUjLbPzkNIUFB3BorZE616IbJy8xjAOa5kBAjf2VuZlZWmWTeu
4GNFM6F8xXaowBME/qBRgNFZBELvqVkhhilDutNv36mnWcIdt/O8YPyb/HSXQvpcGmI/kNW6oTdE
Zbml8Rsf9qL+ecFmLkUcR8Vl3ycUQ3g6GF1hiXtygW1zAnivkyop44oteyURJhLz5ghWjRVEMxVY
SO2Lu0Orz42OOwTrB88hCmZE2fjuYxeyXdylJN/spB+dXgPLAF8beagXyfYgymFOOsoduHv0+rQz
rCnVt+23IR9WlzGw4UbiRDK+uzc/O8hPMjch2AJS3nicr/EMlHdBmVwaX+oSkXwVtID3V2IaMJtd
QyuxcWUlLDdh5F1/KjULJA3sFGOtSGpFvQ3tYAfXbAocDNjJHj+ES9ACBLJMcuMYCWKeqiwSg92N
Y091CHkpqFBgDzsVACelCb4oqgFvcAeHGaoVDkxGKWosTxtaEU+OKhcnlefF5xiZto5J1GRDX+S7
dGUHkBI5kEX5MmEWpxGj7wJj1uCItIEWnw0XJplO6F0ppdehGzPFxrOh6T+R2LJ8YMf8I8O8pwOe
a1h/hU7cA2xqJ0zmU06H46m+KYL6tCxNVYgfenpyBVBwIomyrxySsUwCQJ22A4gin836dFHI1KPn
cfm41x6weMVdI//mtKJ/BQ4e/fy0cRyGuNOLu+xPuMAaYI0ncsf9PUZ2kXK0GuNIr0+j7aFxVqKE
Te+0C8yf3X1Us53kHbd9KM+7u/FwSHFfG6L0VASe1LL2AoeXQ16rg0dQfHFdLNQzCEot4VIkaRw8
v2owRn5MPQX10HTzJNnfx0aB7780pHMo5iAk6KufVQ7P3qD72Z18NXZnCNpBPySMLKzSa9Kld+DF
vg4oUJU3CTcwwsQMUJECxWKjb7fk+HLDHuY04/516CgPGLefjDEXu2HG3+9i52uCBW+1ScQHTjJM
fFpvn2aJllL/tEPBDdxAIVEhIicsY4lNiAawJ4D1fFDvWV0VbZAXUU67wHfr+2izDUbszpSLbLmO
7wpvNtXWZloktnaT82TxS2zJp/dUWIkg754jQzlwF+0+IITnssm87RCeV01ZGuwZbVd15yuS3xGJ
Ipdq1PSIBVbU+bUkXLXJpzrahjGYQh3k2uCnJcBC7X72UETzj6hOGHnaqopTnRRS+qDdzrn0qUiy
h1uXLWCYWI5cBukw47/27Rb62N1yPBBqc5+84w0vVEVXaJXk9DxJ1UrsVeTtEBbn6usoPV/ho4Kf
Gt8hwMa1iW7HYFjor9v0fdjz6+y1BwSzXCdOKrG2VHRbJy8miU/vcZFUFVvuNahUhaoefiGu79MD
KLS+XUrJ6Lwm127hwXVvKCfYWDREC4B0ICQfJrtP88PBlnAg31u7WtVXjiGgQtrIPA/27pMFRFC/
zGFpw0y1EYScknvKY8ZFWZn/UYgu8SpqXgzRwyecNF89xIlCXbTPRWcOBG1RUbABqKTvbds0Nv8L
tDnSFdApYBnPu8XRYZtsjPec1SnZf75xDz0AlyaClBULKQcPWrXdzaIM5XMhNUpNErFpHB391B+1
YS98Rm/VOHK+84cLY4Rr69iISqYEfopW2Rsut3z3r2xgeabQFjF5DJJgRMK1AUCF++Gh2ZXDkBFI
nHziFLiXGp2qWjmoJkF5qMPQk1OS5lbZQls1JlXB9RHX2fTLkugSe7dpq3AwSjBDTPco6ND8PQ3j
X6BinHD9nstj0V3d67o1VnHg55qBN4XLe2YWlDEBoOL3Yn1XdniSpOVVhb+Fy2CgDYz5cZU5eez7
FYQ7X79yyV3wo0gVdrNLKm9ObeKAUhZqxWMnudP+XlJa5TGOIZBqE6HUd+BTMigSWzzOo9FRRhvD
SrSjToLJllQtUKF22trCReZuJlbWEm8XrnJLpUhAWMM7+bTGpg+b9ZflkT2n5K81wJuxMfwB3SuH
HpQ4EuE5Zh0CkdLjMaH5rp6da/K6eshTL3xvo+T9LQPMY8PoZUGE1OQTXvbwIMae1gSJF34rJbFG
ZJNSd7EAYDaLZiFbP0p52EK9CEamoK/WhVNFTsq3q9VrQKbEVpxqVZdaAS/HTTMzBRMUzr9r6CJM
4gJFjm1fZ5Bp6hEcDbO5bAZhK8L0JK5m1tI5mAHmHldNaL251NbBrQRtYmWpgzBPUxy2kU0H6KH5
TO9xrvEbKd6Mm4HzFwNDCA4ldq+RYtDDYspJKJM76JWwIv/QF5FIKLrVZXhRY2MNJzO7RzuoqiOy
SHhAJuZzhiMQ4YIklT30S7vxkT7nr/IQ4v6mojvAqQvQtoPBLgslidBoUE7FpfeoJ8jUhNE+auDN
Rb76IZOS/YVPn+JsVWcZnA5R0bO/otFdywl7Uhc9N1iGlSOHTh69k/Csf0+6FQVcZLQbqHg58i+o
FwWnnK1Ri59LyFurGO8V68koaGEoJy2sjgDJBDoLEKBX2L3tf3lBGyEkFm24RWhmL3TQZiM9jhsz
4ei7k/zzUlJeRIDgB0g86ezZewBv58EigbVvhHBpJ3T0cy89VvuKI3skj1PTytKFyVu4g5Jy1hhi
r/gtjAhma+ytIS8jp8tBEyvBSvvq5vwBKtfoh4ehh1XpM4iERAaM31SDYbNE+nHqOjopN6jNxyfx
6oM64eUavriz55niL9cPpR3ZyRaWnd8oHCla3P/95wswr0aEOpPeDpdIfjwBNQ2aJ261mVTA7p9I
5fztZIAlRZFlr4TIUbfp4MFKQ0NnMxIYMiox+sSC4xoTCMf/SQrHXvPl1UX8q13JizuWVOdBwCk8
3luSe1ppU/I/Q/7j4h0cQ5oNW9Rx1Tev5dLQ0bRzMj9sUtyw7SIv1PgPIpqpNUQMTt1ongatgmQz
vTEjK22HLhriEMwmGC4FGrIFaPPG/QQ3M3DFenthA4qsqq9oq8mGbCfQnX9FUjPFAVEAEeXn4RJx
CaUfB+8LaUNrbkEyht3Efza7+HBTMe8a/9yrqeVt2sPVoZ4h4+P8kYXLVmNNTG1RI33TDmqDMnNn
5d+mt1+UKKnv3Y1yUxupZsdliurP1oUb6dx6YdHuY7Uh2A4UTcOz/8X4nh/ZlFcg14GDFEMEgYDP
Y5kC7CsGJriQKuTh5rGC8KgoKoS2TsSEt8rnhF3Ty5ZfAVlkvfqp+T2K16u3HJxaWlMLuA6rXnnD
8QDkJVS+1JA+0VrBsVUP7VbXxla5TFycRC/GEVahYGmVAzfDHXCOJuxYDpgSpu15k2MqOXyaaR9e
pko4KPevsohuArXKUN+eIQ0FR8v9WYEvTAS22eCe6+7R64GhA9IuJvATl/QrwUceJazrL3FkAKpY
65MpVJGYayeD+5SiEgiUFaHJiTLxJAgxKlKnxSjU54gOZEpL/g794fo2pLX6YE91s03pH/E7RjoG
8AsFGj6meRnTHBSZjRXL0ibHoN1jBkcQiNZ1km+bGZogyupE2uO5Z5If/hECsJOsTpZsitYOIWGJ
gSlajtRIDIJ29gDIPB4fw5S1BYZb74Y/vunOBxlCGHjm6Yl04IrvyGy08zXt8yvy485IkuqGzWaI
l0LwS2VKQ6fX11igEgFU1rzy6Pabw6n1xkjC/ct5G7Vigiidmx1Ed8NfytHzOALd6AFixWEA4cnt
mSTiQ7MAdz6n2w3cZ3xG8MqcDv0N54cQdZoFP1k7GrZoHwAqwXW9Di1rOQx6Cm/j5vd6ZJ81bTOc
bT9Qi2DZHZ8uc7XAayxCPaW2qO9l85zz2uVNZwqf2h6ItlS3c/JEH4g8QJxPYaMoKKroVb8MIkl1
SBG7A74eIdquM0da25v9baubFHRmOCuDq+soqR7Mfm/a2yHvPaaZEIAdBdOpEkmsqssrfRVo+LBp
IQM0vllfvzW0wNjyyK0cB1XCyQWLL8HYczZJlG2VdmNBnnOyjGG0JFi/EEiub69pO/Q2tySTkRRV
G9Y25i+xUrfCQYWvizmagko71fDsHtPbYNoLXMD7LGTh60vCSrTCgXm6yjyJMvWxY+vjfvDJQt+Q
SLQMjtnGfEUSGvi+Coq+aCz2mtWY2SI+cK1uDgdlTBlf6xEPu769k+BM2/1Gy4BU0WBtP++irVVl
GmRd9klqLxXS22e0bWgw0f88v6CFe1pA5gsORt7NyFGgj49az87+LrSAbB340JUF/2HJId/5uSss
Up8TaLyUOkC3A2flUd3I973HCXv7U64fS9BI8obJKAUD51izNAyBPjd8Gw9jfnmQPedgXYz+y5nE
59ydvaLGydJq2/DUmSe1un6v2Cm2/Y2gngDYH46M0I2wGZqtRts8G70nPjQmrqRPOlZGRRTe6k+l
Ji1mUPg3Eut/bFXbY2dNt5Ge3ZElks9NUkNUgQmoQ4oCvRcRO6y1iV7bum+ME1xnIyLYyFa5knJe
/ENYoD4xNfe3Kjva1TPdZjbwhVTONt/dKkDYgg5Leg/gT3apJ7dO6e+5z/A5IDb0JXtVZvRUvnna
0XLj9VR/t92eBj37QfLy19FAZH9m5ixKcVJ+jPv3ZBaJJPOTNKHif/aRV4U40SqDhpArbQzLjejr
d45x3X1hL7wmle7qTSHKBhvk1g2Vfu18kaT5wxsZt5uiQbL0zcvA8dst0ETdW7zgOq12IzQTaQSX
M0306CHYL8tG2no0mT6JqR1US3RQzlLPfuaJJApJ0o25jj/p/laiXMfsyz+t5ToVlVmnHAmwTZWe
ja8Mts206GBPlFIuxbgRfshEZHv9WPk9mSdtZeKkZuJvvog8YtzvrcFvSI5KTaFC2zHBNN6miAYr
DwRSgLm+HES+j6RYpGVQIK1IK/rwD3bSAd4l3H9+FZj/bsBwiqzmgTyJL4Dcc0Vu5q2BMQDM6f6C
8BcNw4JMexdlUSez4+aQ1QLMeShz3hd+vIkMJiN8tPOJ38g+HoOGpPmIUMHnprckQyDO9UXgYwn/
mRGgIVPbiaT6nxfCgs6/gZAUI1Cw0YE8iqDMc/SSfOanPjnzQGT7caQeucIUudPlWer4wqzp4JuO
wwsIGlqpFOJLwLraKCu9eg36WpjfbgxIUFXkrFPk84Fuft54SMmt7GgO/k5bU1juvzH3PRGHPwLH
/SfjA1ObbRGF4MuW9jDkbMb1KU+HPkqzto8Md7mgsyz3HLBagwq8grndcHBSmchLDZlkJ0D8a/oO
+2r+hNpjTY19XCLFBAXNcCSTCUsIeioDvRaOVoCvG8MJ9xlG2Vm1AUBaefgi14frQtvgB8EEGgBU
rQVjDmW2eOCmMsaA6RsyWHC1L1UViMMSQ+TGzgYGKe3xOgZTqHdb9gWMuVqqvS3ECaQsVOlcTrEb
LDqCX82Enfd4+5nyN4gC0XWkbSfuDxjI+GeCxSUSGQ0gEPts7bFfvG+Azi0YFTxstOoCfyR8lGUh
cwpHglq1h0rPgy2RD3Nd+ZGXehXNNBDILSgPYPwo/JVs09Qtc/HSopP3rKc2KwZZlH63cEqF516Y
YjDKwbX/d+iG+qvyYx0xSE4mTu6K/+qNxlObn0cemUOMXYpr2fT9yJC0bxqQWzAuRC5nvZbpgt2Q
lGssWUvcNyn+Q7NfUH4WXDOYgbAMysrO43vCLm3B5ZhX0Uz8gorpxoZrk1TRYIHvgrxJqJrDNIJ2
az6QAmym6ScGUE4Ytcj3Pm43xXfnU/wjoWCG2HbjTl8o2C0vj9RNssclWrjJNyPgsblX98CHhPmb
ujkR47jWRMf0Xfd/zxeWfwq2O1gvH+M6NH84fVR/3C716yaiugmJ0wMNNgxG4JY9/ciF7hd0Z39k
m6KpZMtRvn9PSxz1msTeQu50fR/Pvog5eup6Zvo/Y3/ukctMaULJaOi50CN2LbmWA/jIoBTLObPY
/WfxOWAs9k85PB1Agie6jrALILZE3daextXxCJN45FJMYZtXCIHCQ3M4+OV5k3P+lW8Jwump8j+Y
9a8C9FyB0JWKWXNEHkc8zVuxuvjMRgShwGmql5DCUzcKQboFUOyADzhFW2FTipcU/C5JToKvBRbD
C4wVD+gCLjRdWyx3tz6u+BI2y9a5/YS4wB5jgXH1BVtt2Dy2Fi7SjzvRibEy0ozNGgVEAmEf29De
bkeKEPzS9TTdfOIv2qKaDoLxoTHXE0AHsR0Cbx/FG8QOiS/tr0QYoEPHE3IxfIBETr07W7t1Xh8Z
HErS71nDu2Ga4/EZZ2GCtVjQe7hKSqsTELuZKBJlV9IPYelu730BEqiauZlyyrCSJGgcEJgGNEDy
qjWK6GW4/Bqv70H/ZKEfObOWT1U5w5Ry/LknEaDIKejw1AFGu2spnW2EVwdsvjwE/2kt4wIxSVZK
KgE+/sptDXO7EtSea0Clyf6Leh3iXcsO8dJJo9wfuj28BA9J1KdDoATksF6XVzOjQneCS+bz3SGN
ghjB4liNQbok0vKm6GEhtO2UNOwcIFJx7UUBkJC0Na+E+ZmkaUM4jGRDg7QoKBat4pozE7NetfzR
OksuojGlr4+c5xrnCrZB1+840xw//yYocrLX6toDJvxsLc9W/xHXzwgDi68ekfWAnmztXum+xuLF
M02NXIzG6ziuVrNrvEM0LM5RZ32ZmBIKRrQt7akqSyymlEZILi5MmRz6QIOAwEQhb34hE9dqU54p
oHr0CNlo4Bnm5sCbmmXY4iCwz4qon22PgXtAgnplP8AHygPl8YFYe4U9+SObPdMiXdmuxpD7vqBl
L81L5kbO17OBjpFla6SYsFmgt83MZLF2GyXgsqta1OUETzDOJTVf8v33bH7orP5YnfOZ5JgVu3BG
bb9pSDuF9QIzOXPCQvZ2v/sFCJ0z5hZ1FtuXsRQDKyy1j/MK9H6nbPd5DDwW23BanDnqgOePLV6U
yGqmN4B7LHoSfOBIxBCcP646s8WSD0ZBVarx8FyU31tj7xPY9ppfrqipMsYw6HRc1k5IqFW4Dzpn
93P61n+42F8jvKhe+L2l9agTkvtExAmKWirP5hrCv/gmB8bApUEbVwJSf7xZg2VPJjJskf0olTgB
WEI5GUxI9B5o/Wbxp7QkIvb3qeOOFDyBrTMeZ7DuP3Qx1rgkgusOOSPYI2B8llDpBV0FdcdbDG8x
RuY5iD7KwQIG93Roze075oGPKhPQt8j6Fsr3ez/KIpKGAJbiZVZGzjO48I5uAHlI9j/qkHh3qebC
oW0F6rj1zDFvzVtitZHcJ0oaFE2g5dpdCzt9r9KSM90yNAQPfZLAuKk1l89n8gr05WhiMryY729k
T/uqk9mM6hCgDIEweoAgt6LSbYAcHb1x6KIxMNNrYkqSk5CK2Aif8/svVduI7hHsiaSHYhRH00Aw
S5ixFhCOdWzWxo0wo8vIAj62e+mlgQPbhHF8pykVBLI60KGfH48MolkkkJocuc9OYIVLSmf5rafH
+/y2RP5vBscOMlwUq2tzU96R7/Pwdr0dgAKtel0TYLDnDS5794kDwt0ffCVbsKFn5y1jH3r2nPbG
48y8dq798USIjSiZPmW8xzDw70ycoN86mt0en46pt3HNye0xUV0OHMVG9V6+d2jiGJIc5Ptu6Nyl
LPpKkhQlW8+pE96kCTkV4bN1yWjTa9dsw53gXrFBocf4u0oeoB8PzD0NKdo6Bjkh7hsIOCvqv4Mq
DDBClCi2+JzWPQLH5JdS5pjt0G8y/fT/2rHyD1c1t5FKXHiPK0wM9wiGGFF7KFni7xbzL3Hbl0yh
NT3fmO2/tPcsJiHW1jCjUHYdssXAsn2zlue2LjG+eraswhpe0ieF/ZEMZ+QyhSLdKLhwKAYfRFND
LtoI74vtidV3OSaElX+wSae+naVgUxt0FhU0zxKJuqOZXUo8bVnsOxXlJI6XNXSGp0HOKHxg0GId
aFHVXf3VU9P0otKKDFcS7+ePPoEyhLTvcSFAQNKJZgMi1luHQmAwIqi01Xc0QtyQAeYCGPdCX+8j
mw5LkkmTd4PQZOIP63GvFJdbdaCz9INNBd1Wlta9kx8Fs+TueCw8/poRrgXEBrZFzm68/1VipPOV
UDciNXVcOhA5GayQSq8xv2gcZ5tabXm/DkY7IQv25Qf69PQJcosg7KKTsw63CKQ0JFLhIui7i1Vl
Hf0duFO6INjUOP8hDkVmsC0m3gmcySUrwy5AGU6SI35k0Daj0GGi3N907WODpvGrxXP1kAGOF/G6
YNOh2c3+CY4kdTEeg0ZZQ/zcqbTuiQaq2fk1kuijTG4fedSZWxkUFn8ZvA4Vb+BP+icJzZej9HZd
FopAeu/Uy30cWwchjMxWY7u0QmhMpGnuwRbh+A+KlZDpHT7SgbjYqShyrBMCYoQHlPr98kZhE9Kh
/oY/eX6RUdrqCwCZ0RxCXtRb3F5sT9Zz9VEuzT+ILDG4oC/PPFVAugxFadOP5921Ad1YxJxUFGmR
Wf3C/PJJ40II9GOfR71bZOI/p1vRNW810RHFvBvdLisxbgu7lYp1vS6M+zk2166Z7+lxVpROVAX4
lEKo0RExg5cfUGi6i1yRp2XD4W3Uf/lOOV3sLREfY7vl1G/6ecrjxyimWYfbOJDEU3VZOkvd0K33
ZmFmu5fX32FFNjJ67t5W0Y3vNBdQYP91X/2mCQcfkp0V7o8p0BNKvlNaBdRtRze0RbRYsgX+VZi6
Y+QxhMF86iumMg6eajsRBO8eyLlQt3pc/3Rnh3r2I8dwxWozdW1XEBi19IvK44hIi3LA5R2Cyu2E
9vG5hZCUTcVnfhebxMB4cZfR6iXM0lfoWRbVkTJVnYzJ2uNOi8J6iVf2gxQdk0jXQmfCmMS6+NOL
jgxEUG3xK/P3G4ekwHM+GaFvW/IDooxBVPjO4FwUJPLN++crj0xoBfALGSmRLFiHEkoCEVXt+bnn
0WDHYikGoNMxPZA08kc8uNT97Gi5yo1zQFo49FjURf/xyIHFerW8naoAH6x0OqBPfx6Oo+v+F4MX
ra+uMGM3Kz6w7Qu4fhsdCo9gxunqXpuzJNEQhoaB+5ecI/g/WAwZS3XB4uPFrNzYqLhygTBiBIjF
mMeTMU4jyIRPK5VV5JoGNoj7a9Ci+8gOsg4mg/+bX29b7oJSFbuMK8J/9CDzH2UWAcEbR3WiJode
Es/viwbjQr3zkLB1PmQL+bjv7satWxrHeWtXHF/gjNoLBIzwqawPFO2wOr/a7luAN6chzKXFdmtH
Tn6aVD17w930ep5USdRG2J0WIYDGAjl+EfHKKDZt3aN3vvi7KUksi/FpC6mkLYFHE+PxuNmaBnaY
5a/401bb3vU4ZnRLapnw7EffIXZIcObvNpH8hqyelffXRY111X7/7sdfnMYnNegGksISIsJWEPt3
/+VfwQi2U5xxmky5K/RS+i6d8Bm94lQrKni0q/5IEvlPOKmLFO76edjgxhowNTvHRlI04jtc/8Em
GIabCXbMbgWq9jTZ/+8jP5VHQF184nKj+kz0UJT+mAY3qXVMqPbspz1ptpB5/O7evWGXsmdLnRAC
k1ubdHIvP9ehO8UBQXYCXTB//y1o51FuAAaA/ypEw0vh8Mbco20ZT1OizQhmyUu7X3GQp9DYR2ir
a0F+8CpvQ2p+fFzP7k7pWnbW0gp07crs2uzJBdnjsVCtN950U5iW++jrbDGiO6SszklAPIc0KXhx
5uGOVBrbNDWkBH3g7a6AZnB0zo22s/oSIWUGr1u9JAqhbSkdF+MSpJnj9WqrKNlTYfJfagd8h8e3
Gap619cbwTOHjGuPEi0IbazpIYUS858/a5t7IyA8Z7HpDcD/oCTTHoiaGEWsRBmOblfZWJRdNjnb
JjPbGG1YIXHRSTvJP9rVFvC/TSBX+//Qhowl6XKgU6VEjsVnFhJGQqcSMnmWkn95ZmcGUjzSa2df
cM+Ks20m4BlCqwYumThh39VYaoNXQL41+WHKag8E+1im9a4PbGhhXhhoBAVJD2aY3oupBRvhNJBa
vawHPEi7L/H7+Hir0ap+8RsDGwPYZkLG6na8cW5ac5zYetIkYMSEdc2InFiT/luhl7nBEsYXcUJD
q9wfT/hReHUiGhDI7kqXIoPV+RSY73IWAT/X03XZasVQ2mSRu0FEuQLZkihFSJz3JdFBIz81n+wz
ETiQNGqCcfFejqC+f6qNQcuTNGh0eAMSSfRKPyjfhEXCDRRuPKWtIxWAbCdFvkNKopa8YVdJb0Zd
9vt5mKkkF/Oq6/PspvmF7T3b53MoIJA4hloVtN281wI/2zDlpdMPHR4VnwPD/udUO2a85WtYxfEA
e9y1Yl3gRO7ghTLaRBDZdNQTZ0Vj7nQSlAdYwvntHBTEaVx3EWAeFPFThTlSpYoScwx4Pb6Xqnzc
RvwzkJ83ucTnHI5oKS1fM1aPOrs7Dg52k5cchScSxEhxbPMUlHW2ZcLkxtkp8x9mXqtCNMqdfJqZ
hSFId7/4uljYRJhP8lvCOygbS8fGZt/5peIzYpuZPUZlMUpCevogIcKySorse/uhGNryvPPjuZR9
5ZF4c69x6kfWHUKBb6wjNd89vakZ7vj3smCnQRz3+aV0N8br7expTb4osJjuUeOulwUodUoOlgzr
PVjJ/w7qxptp+xUZJIh8psPJnWXnZGZTszi5WKiKglYGg02bJHA9tuBsSakMydpmX2fBXkpM0hgU
uXhTr1WJZJaczqOquqUmQFgQ/EkghNUKyvmZYhHjC2+HqA9S0MgDPp85jcJpzMorCv8A3sjNCmly
Hwt5cdQEd/NNr0RJJxofKTGHncsQi75FCdEPAM/JUdeCbcUOyf6f6BeAV2fH60cCHgeIH4LlAvfk
98KzbcUWHC7j0RpEHPQVGvp6EvRI3piItvH8sdbKr50fISep3+GUYZ144iDCt84LqsnQTxKyss4+
KMomPSMjCobXiQYq3XvODfALrpAqruqM+/Va+hj41aR78ut3nIWXZAhngkI4MxbtQ3s3a7ckqK5p
5pvXVO7x37hRYaqwgHaPBfwe0C3xkhDObRf/KwZPSkk4xxUZLiZNJVIF5GDsOM/9T1NO8WQ4wlFz
w3G8yAl4KDFBVfLNP2htrkGYVVGVVTbLKq6oV1aY8qHpvN2Ji/OyTdJ8pa8zO1GF9q9KHvcsSpw6
cxPHpEnDCXrnC1bD4h4zXRg8PBX0YetACQIjgsoxx30N/vFfgsBSBU4PZV8lRzAnYDB+IEdpY00I
rpg/+DlIGrudUUnUCjq71cd9Z0KLadxpOiCXYwoEYu04k6c59c6WezJTa6csRjiKqF6M0b5rwWrm
PjyONmx9xcA1XPWMF7UP3DrbqzwCcj29bJE3IbXovO35W3/YNf9bSi8zfRUa2dWjtNlpqF7KwV7k
kD9q+Gfg++YkiU7VyO7v3rUi4q/ZA/iq2QOpIy3bbTCaVBGI01Rk/fdtowEHEWSCpVtFEjd1TtgH
UPjSJJbsfpwJvCeejzzRLhnlEvof8Jv0xRIU8RDyV5ERuizjBykhsB7MUmb8At2hGAckS4gzvJkS
xDER5JqnxEbniczsuZKczphJex4yd+F6KzRaqTd8G+ZV/fIQffRKpW8G0R4yjCkz9rWWTsIRnP5X
DM5reWAhGKRf5JZHj0kochHp46M0oFyPPqnFwN+lE/dFVBs3bgFWbws/fjirkkDY0bz3C2tUgI8I
yzjYlJpliQqqNgbSHMFYl6k4LetvXEi1j8+J+D50yGOOogHnsHuH6K4OL7N9E1dOQ0GXQiHLjqZk
e7vTc4VW1GVcc90Gl20SLTzjOMB3jGCPC90yWTvmF9fTIywcOg+vWHjenfKlpu6JxiP8y5llDP0Y
z4nd0E/xdibnNds4tyQv5upW0uJCFVkSYuipaosByIyO4G7uN7kmAjM3b63jpakSXDBfiAT7Y/By
q716Z6SeCY9J7XSu7Af3qh6PEpnHsa+0FWMIK68nYn7oMXQsb9vLnZBUWUHTqEI+ltKQ9wPD4Cre
jahY4V483wiisgJv9RvLp560I9MYPTfAfy68CFmS1XItwczSuz4tbwOXOngxcZ+NidB8se10k9x7
HGnbg6QsMqHp1Z3bk+SXwe8FtQ77FQctfYSUBD7tn6aOYem/J601Z0bWP1KMGWD9MCVaDxy8r2d0
uk1aZMa5hqdcmMBWRKjkMxABxaInKpC5PDIVbJ+wkdimJ75GWRudp2WOY0vO/6jSto50MY5ShaD3
Yprq/SfW2iRc7sQaKWm2MmUppFYCxcNrKd9J6o7JEzvw+5K4E7JrGC786RLFBLSEtT7dvH6iz14W
DCBFVr9ot+s0wme/qOBBW3wOyHwYbJgOCj5WpkQf28o2ZM7OJQ1liP8Th74+AN4/8OicG9ear7Tz
WHiAqsZNq9ZGu5UclA0C4i7Mur4DrboyUnp8Xcd6GFo9T981kf9VyhUoD5xYPIZ4a+23vjmgBC1R
pizCP7W3HmBwZACH7NAwMLfcMoc1pK+B2Q9plyN4kOUCHITyocDlh/qy2hbHivWkm8qKaZ0Hdo5A
cuGxkV4PJblxmbGpA1fb1SxDnfVKp4C/a5QL1uivyONcvUlLtmoKnlx1pQ733dZHRz72oTz9EfA6
NVN1t+jiT9CG/RHy0QtnOgB5+wHc0UNyqtx24HiZ26BfMnnJH2t9WvWbK9QRoNoDdfeJXxYh1+dV
8EIzzVo0m6EtiZW/FUyyTnIJuxSHk8StaNpCY7AYLYYjFEBSySb2qL71awSyIRLfyE4taH5evdAZ
xfc1OxCC9XJ8y5P69qyaBcJBvy/BqD2IO8ynwVrh3SHTPb2hR+Xh9MiZFPgHSnV+Ly2+WzYW1ZLt
3FZpa0OM3A6wZEsFG0f6oPKz7eYkRvl9ZMdl25w480bo5pGvd/+CYUbDmQ5OiBp2JbUXfCErY8mI
hd6OnfTqwkVV/YQVii03X74FElpZDQEcEcSMKntlsQc4NLKase/lGVMLpJP4bHfxfzqSY772JqYF
krGd3ayV8l+oL9f3TF4TFwtBfjABLgkLNuTPYvpmRyxApjx/zmjWK1p9lgtiGvbW8y65HBa5d8gU
77kgkJ9SvbUwguxmwL3GtA+9izcydilP4LYFRdIXmwn+NSq62BmI68HyoNyn8ogH8AAerC9x2Phy
CTq/SrhFzztrQvGDrL4yO0xg3pr60bu/+UyQ+GO+pEnMK+4WD0PtX2akd3dGWM2tvqnZSRynCJXY
eNF1J+8+m25uQ79TLws7cUKZ867hliUuQTOV1fBfudvpXH5fZVL+BIJ3aOXKpHBiCHc4SbBNIChG
SYpaVR+mnzeX2hVzKVWHQRiTS6DTOv8TKBCraMr2P+vsn6WuuNcG0kC/uyo2nKVH9nxEbHclEj7l
X9qnhVP5XqJFUpn2StBFCo6hBvmV7PFmUPhHHToWtbia6qo386dxS+aulYPfkRdGFn1hhqbUH6Vr
d2dU75XjthN1t/oUNc5U5VPfxVaZiOo/mNBCPU/yeNYUv78BwGlFOLRMzXKnMZzFHtUlq2SVbEjh
AdtU6TkltvBup+04DoxdZ9o8w4SI0d0Y0cdggltJHXGqzVxxW2LCIoHVOoJjydD/eymOtK47DIsI
Sp6XIza8bQTiUUqm7EDk9zQogSbs9dce7yaA8NughwJQYCDCnGOiyHbvpiPNBR/G3O4+g5O8h2hI
qXeXsT59CMWUqQe/JnvrKCrqKsPlOITJfg6PQdSRciObAs6QWWgMSr3Vtxo9guTar4vOCwEuWTpO
PZwAgPoTUcob/kJ65DGgqJSebdUwGN+jumhtUOuGfXLaZitQFjREVcbF4L/rMQO193VW1F1klXWD
VJmZUi+Xqa6xm1kEbuF11tQiOw+J1TEm7q9KOl3/kBUwm8JDHAbG843c9JYS4J3htjCGquz5F2Wm
MLbA9JvoU6vH5l8aTokg2AqzsF6FVjesah+5pdJANLKxfTuPwbbKdW/g4LHqoAZqxYk/n1Jrzx1i
8En4PPwCvBghLeNPxTSmxSY6DOcWwA2ZN8fXZr2Lxb7C3/3fXZj8TQV7yrRe6nUcqhEl/tSj+wNI
IkE38us/Wn+UN71FgVBpM+0uPBaqty/cTaZm/+zRV0P9u3AuAA2OvKt4AZlsoZrWGoEDV8wOqwFY
UD4nPj5nKo/YW0xgNA4W6Qv+SAOp+hW8YBnBgClo+Td2xOi/P1IrT8mNY7CB9WFl3YE02H+qRmkt
qkuvrS+Y/1NbgzO3X/kZxIU2WgW86IvqS0yCdgBm1AP0IIH5xLxm7ofO8MmBgHctexYConBvK34N
u5RFss1Spl+4lF7ArGZoPRNgyQF23nUvhbY2mU5JMDg9Tg7B5brb6X5kH3IShxd4AnEdEdy7CW2r
vqNI+ae2RbXrolh0/OYVYwz2mwMfD6aIhtLOk3Hdt8nsawwBYriid2OXr5p/Yp28oZGV5jJGUVMd
sF4dgeH3HS2I2n8z0YNPidryuqtx3EMAAjnQ9ih1DoqwrrOXjLTzOS+vCdNbpralaz3G+jFAqsrf
DUr1TMEZH6Z9iXeT46zja03uMo1dYW6N0XUeekPM1o2fVK2NocXSbEWcDSv+f0JykJ+RW45o77wJ
ypNGoHWsTRNXABReWBus0HoPjJLoTgqOcwc+DtIUwyLxkhLlmmtSscuhaCHLhROfbdk5hgX0Szoi
zHLC5L8pAsW18csF2UehWEgJIGIZg5l0sVc5WCt3q8rfMjzmsYnS5gZlumUg+hgz2/AHGfI8DWbr
YYdQEzQwtlhuquoVnY0wPpvR/s6MLL2/J01l01azYVNGBCEvlGAPCCwa2iDJ5H+86Lg8N60tMYEo
QF2kk+K+955cJ+i0LQcUg+gH4cZczxWC5SBeM3DaxwYtPlu/v/bdmyiJLNS8FEj7C87j/qu0UiiJ
0uiPuOfYzrPsj+iE4eThq5xUZgQkyF69YRJExhgvce9c7hqQ6gnojaNPi0l3GS/GnVo9jS8M1e4A
m5oX6DFsh2y6U9p56MKGNq+n/v509fk2w01vjo6qj3UlxooXfGWBnfYtZ1DP6MQNrVadoTIWTHqV
OCw7a1wBmuV78WLV0F9RbZpVYozj9ScU/Wo1lseMQaTGoG71VF2rEinmpsNrCFmOWy5G1pWoUcpo
JR92VQZFI1crk+U8B/34RFP07U2AT4qRm/TNhyRKMUYxg7o7HYbYd+gkc2Dmhoy8liYXsIFpeJXS
HESN8mqklo3lXGYFHu7JPkFp+XXdH09e8MVzkCZTZP+D7b0ec7FwSQ5kMaKR/ILtNmNfz8p21TGg
6CeFX7/v60Pb8tizQcWcQhYQRmh3jyBNeXK3oHYl7017x4co2hJX4Lp6zjCfP+bwyl433zLFFmN/
f0HK2uu30MNqng1pUcNUpYZE2TQOo3tw3VjIf1/8eB3gcAVTskJKTm+l1FXu3tjzgWwdcdZW+VoK
Ad8XfhiIdmcxx/eSSpGWnSeKf4g4wPFawRsMjLGcO+tGCoAgkNhUjgKmlO8xuITE9DCbAmJEp+C5
acSmgDs3EHOqZTQb3xDvfI/CSC19eZvUNtDPgG+LisHrbz3NWWKq569mnMnLHGtF6IQpH+QQQMBI
5RZQq5sZ0/UVPnnyXSixEvHVXRMvrTtnwNuuN8O8+EHijO/3L+UsAJpOBpXZOpdQw471tnGriElu
lVQrvpN94xM+HwBjbV+HQjB9UVg+UK1c1OmYR2X+4SSxY23w5IxsAhj+F3SjTpDuIfrz7wwjkd5I
mUqR8BaqQCmezUVnhiNXWhnht2VMUbB6N22tT/G3XU00XhNMkMP8tZgscBC4yGDnn1pu0Vc7cntz
xHWKSuSLyuXM1/yToyafvOye2WStr9LOV7uMTpZv0SJgL0Tso1W6WzMZl7/zybMTKPYLZEigonkH
MWgEmiBKbdDIW3P/CgO1DF0NGs02WQsLmvwz7fKtkiIS8fXVKPfhdlC1/TIwoDBqKR2h6oEzc3xP
oxwzd/DQdFl9G6f6TT//UCQsswtR70+DeCqYOsnBu9MtDP9eFRDgi9VJGGkv2yfXG6n7z6IpOIUi
0VVldtPEfuChJRPJkpHgTHB6djE1Q4SkQAMSf3Z1g/XHIB+dxahaMf7ET/MnRfloOeqHywJiloUC
IoDngWXijO4OxnFxkrf1qHlOb5K4sffmYOTWdNSs5EQNzydLb4PGvGZEw7ZYbw3MrL75wXEIdNe1
1bupOOFhELr6vfVuS0egfE8cO3/x73A5LpyPLeaChmznkljsj+zKXaqcg0t71jCKtKicdonDpKuD
MrTQklrt06OqQCtHR3/ptZo4TT7QcJlVS4TlBsiQ6QjDtVaD6Q2Eq4pIjTgz3bi9QaP3ZQOACPOj
iBgtJKjlrRaLi4NvEywUCtdgv9Za2arH7x+iBr2J65mQ1IULq5hQT1f5Q6v7/lgeY3eoEJmLcZZ1
jxD6L/Dluj1bLZLbWezzrH++m9J3vd/B+tLYcsFyUKpzSJAou1nT86XCrZUouzP6QmgT7dQcXowl
ihi+I18Ky498JdrC+qqNGiZ5wYIJLYl5RVmzefs60wyGEjGbpjdC7jwkxYgbrEo/pjXKfviqGvGA
gLxuxiUt9jz2/znCYUcz5T3Ddw3ZoW8948ue0+bXulrcerethUf49D0wgB87RJX/fLWGvh9W74+0
MqEKWELtkCEpWNcCAXeT40dzT/gVIr1Xev4ZUd9qNsj+upnvetbDOw1rZ3EOJqkR3JSuC8PEt4wL
uRJma+fxhCraTMlCuPlkGd6CsoN4tbSDu1RT08TpvzeKN0ori2BUl0axz7tFWYU17gf9ZHUlJiJe
1SQ+S/b9nU5TgG70+AY2J31nzLb8EppbV24s4JhZFR4dv4qXQR7aUaaenQP9drzLN03SUKnLAUEm
NtbEaj6nFaOcWIc/ADkbkXpDqEqi4XPei/Zc2nXmFVi/WLoL5xcy4ZTy5mxlG+BkilLSrKWer8KU
mSxc1PkVLMInQztVcrdKaVFHfsq2gaxcyiMCeLzM9Cqe/5MkNMrTli+GnFziBVqTp0XPFABXHwGy
Gd4iGZeP0pNAY9ToNqwRl1fZLK+7oqRjlYzBU4XTonF5pASqYGX7CvMBJcjpy/rR0ftElYiEf2eC
U2qw/4Dd2bz5MXBaZSayn5tDLbMlypyTJ6zDz7tntVO2/Z7YJcTW1kV/ve0tb4hapeWhl5FElRFP
g+UkX6h/vNYnvAJrKgCAT2WCcuSLPz0RNyfRQkhacft8LIDrUJMSpj5/vMhwK02dnTQ6C4hXqwxL
D93gZ2wPUS4S28iYyVRwn/yaVelLpsqCCv1kW4Ug2I/Ssa1/I0rUHOTo/kOxvutMHwuElkgp7DlG
+K1cZpOqwd2XCQJwtNM3SZSB/MsniDyPIg0HuU0hxZUwwGDdW1rtZSmVJv3dC85vXdEzvQ88xAvn
tbUtjbzMXVgd/XV1oN2+S5fflXBDcd0AENIGdnsfQEap3Hi1SmJMmvEloQbvubkamngZpr9p/PLZ
3GlOzP8iZyb9yo9UQdxIg9VKSPaiuuQVI6cjKhUWwAHSWTAsJnt/uPPIKwqWhRmgLeAUC++EwxI2
AIitvlJlhEXXqeuNtta4iccdwoCWyAbdMNGYVVLk1gt6j/Jy2YaFwlbBbgJ7Hkdg6eoi5cY6SGdC
aX0d7QJX7K4Z64DJXHs7V55Eu8SFFAPj5m34bQJK2OtG0lukSha5OXaIShAUuMZdkPt7G3iZ/1hp
baH+OEZhmu6/e19bfB+BRzA7a+1jao0o0hk5JGBKXEnZfSeLOrhFvG74KN8Kad7Qcv9/FL7uMkMx
VwEQziDKLL5fGqRg1kNM/LnyQRDe2+w1Yc3sBIi7tQuLm+Tqj9yNgvyTiGJIAG98h9/XR/SPGsp8
4nNeWhykhetAEfr45P31gghz+uyzk1Hwif8IPm2KPmNpFc8lp6v65VyoOjiz6mqpQmFrB9i/Cbs8
1A2dpRf2+9alIGMZH01J4mVbE0Kfhx9OBLYLmt6FPp9sPCBeDwEgTxvofkL3zm1JQllZiBg8inkm
MZWj3hmnUNqfs9+ND6Y9HuyyEtEl4axB/UlPpRScOdcbclYUUz869osd6e0m+1mAxpolw/y/d6vE
5MjaXqENLHxALqurNeXDn1oMSssroHHVkAUedY+v55VEqtRQ0xxcyvCM1ddxZdN39kQQYbqLZ5bo
ZLlEcCMa95I+Jbn7mKfIF8abI0+fbgmYmaoOn9tsfNqLGTd1l4JjzwVhDDDnAmkKU2/wkd9jmr4s
1GwcmUS/4R4bQQQido6ZSgljPNLKGgqLDIwEMk9J4kW7JGak9yQzaav6wOQvZCqgSCbOam7s0VQm
J3keJaMJ+PHkJAn3eU3TGxZPdumdrwEYSkZ/fbnjynHXfjkaL4hoIfx3mvCn/us/D38uFor7e87x
QaIBWqxagoebCBQqMBWSbBxJdEm7epSKWbfhqtJRaCvJjXW0csRC9/2qD2d0Htb6P/Lqmi8uQZLZ
UMnuUxuXfhI3syubT6ady6CwP92wE4S3573iHiTopSzOWJJDcUcvaeioDybVWzYvRHPrG43Cp7/b
FUTUggj3FaBNrRdKJLkEmrzf3+TRPxWoy5GskP6Xa90tf4TcZtxfUevVkv3eBsLLBdKpwAkImoo1
Lpa59R6XJ6vOdmQYMrmUfHBRecSy/uaFOsdU+ix9BZpCtfBaO7vEWbfo7QP5bcKT6zttbi18lm44
z+m4eVSGhaYhD/RJk6vMFZx08WZq8YuLdFwOGm7jji6Rr99rbCkLja5ohen1gMy3vCDIWTJzl0Da
3no5MUU0P/LJZx7bWb5/HxtQ324rZQ1v9+3u6SuKaL31qO5RHJVsPn0kpsnTT63D5RXohty6Ee2k
2Bnhk33AisaQ7DMogD/9xrYyziOq37BuTO6QUIOz/eZ3B/g6teWI/8ySq2LgKRwzUNebu7U2xWxj
sHyaTRWpkWbO2XDiX2aRWgt9vlL1FcuZzC9R1ny54YlYjm5EfLOUQxBst2rsoS48zWKK2MR1StUL
N45WKxDNd2DyPLV2M4SbsGej++iUc7ETIkl9m8BzdOOBioRg91nMBV9QeELQ7gfKABol2ebdRjwb
HFGXAcaw9ulvYVvy5EBxXNrPgz+LZnmyQiJ7iHN6QFNUBNH2zRkJ9r9nXBQ98l2MU3mRgvEb79DY
vcPIsZ/BFASzfhFzpMpDjOibkCTBDLRyimit6MtF8BtHyABhtLuZeH7IfU3AXVdepDDWIBA4uhW3
uKDk3gSWLIsj/W8aHasKr18LmZA1FHmHGs72nH1halRgqHODDWNnGELf30JM1Wv8gUHL1NSNUiXT
g0JuLWLeSSs90RRj+tnJ6DFH4fqV45OjbkNKjryWLbOkVP6YktQ/llCx6dbKEyuYIvUX/pXy5idP
U7RxVU/KpU5zP5VzQADdGQvj7ybNU0GpKWMoYy9MJN/QVEwNqbkWvPIcL3UymKuCghBr/6Gh1HMw
JvnbozCOhHAvt4oA9TbrQnXZMCoytegGIPovgnEpbUozKbC3wJJ+ee8v39l0xw==
`protect end_protected

