

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dtD3GNErsQQckBQO5gsI3QX6KEV5E7ts5EyKqLUcTl1nwscBhbrWkPvqYWMRydPjnBTBoa9evUwI
eW27Fq+haQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oFqCFRLETxY+F99DAnFXOEG0LNv8AH/BR3YZ6PVXco8GYLMMd9KV6vIm5+C+Vn5HY+mO8D+YQphM
iT6ggoff3RcuaQWL9i3ZjDl1GBRsEk0uLTUs9Kqo/a2mHug66MVP4F57SXjq5TzXcKSiCGzszvr4
UvcN0RMZ9JMmnhPbL88=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dUuCsN7w2Ia7j7Q0zaUBQsXxD8yReQ64sMeg0RFnfoygLxvK7nNNhyyZ5VM7b2BhPDex3Y1+/HUI
RdTBcuNkIHefWDCgutTO9TVEdfBY0xOiy4OGbsX/OPTDnAl0LFJ+EeKTP2u1KI+sPxuNMOr6ZAUE
xOxk04Yfz4CZB6x2gMQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xhN6lxizkULPoPRd+P+1Jgxd43aCEBEjYwquDYSQqwPtbmDQoUYoUVKq7Ucgv1UXB7oXSEDiOK5k
UiRNNR4/JdOEYKKFMdbk+2DdFKIt8zvOj6Vy084Z/twNrqcJnvzNIyLxBEsfbYcGK9Nu4QmNiP5j
ewWJ6sf98qt5NqMv30tVy+RX+v8wrK7L63yG3hqyL9j4Q+n9lfxzSTQQIGHS+SYp0NN/+K2/PJT0
uIubVtrxnl2QUS31aKTOVDtqsjeAaGsM0OZVNqDXuWer80fVF7Q8zBgYfEIrXXV/13MSal+q5q4v
wJJfhAhOrW7m+6EFwKbcAXNla3LO2uO5AuXj9w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
riDHupA7EDOiidnqinxH1xY1/c3WAySU7Hh9YnDukuwyIlGMRngvANBJFw+wbARkxNJ5Mop3eBX5
iC9q+75362b91X9QGjDpZjxLCuVZis3zLqDK52AY2Rly6BKO5HoKAmvXIUEYzzWRMNi1b4qsQZR2
vH3GMNcnvFUhGmXsxSKsG1Ypb7JZqfuDSsjRlBY8VRvCq1BidT2PBx0omBFnNJb1jqKV1rgDVQfK
IDms3jRfQKzBFQYQ74G38cWYQHO1b1rDZirv5v+iB+z0ozneNUYQG7v0rP2uDNG1uiPCFKlDisFR
ncYcLkKyw9dVdzITaPdZHnG3mUAmDedAbKkzhQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E3BMI5Y0R9sdenj86S41gekYAgvOsWUAwBPXMQM2N9bjHn3fHL196RqOaI2vL0OROC/MuGIrq9Xv
vUmCL/boBG9zWccOsrwfp4FijlBojaTmrgC2ziJ+2BzXT43evs+NNB9UbTLUKpx/JTajjMvPa1Lb
Fn3HjiraVE1jWaIccJRsLmB+e9+GuqFZ2tyIsmgCO6Qhp9zUTAWQNT9hX0+OCLU+BjTug+KgDkAt
gbIHzAKcRjh6LG24DQm3ZxQ6cc9XJYXyrx/MxQ0bLVIzih7+IWUHEAXXgVtxO3knw0LSKMNDPn/j
iQ8C2+790TlGBlZ12ewscMR4vwYGvY5t3HPBVA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504720)
`protect data_block
Pzj8kKA1g9GIoeqytZobxLDZRWGcJYXADSLo3ud10PDAi5NkJsDPqFt25s8uYVJvpU2kFaEJsSHr
/Q7uxF2mSPk2WUmKUj/0+nSxCDfjmPsfs9yzrY8HX7GgcqsvrznrrflWelnXFSlf3iA5Mab6ZadA
/XeSJodK46NEwLnuRz0ejPvWAg5w1lnfCviESgq3TAZmn1QvzN1jwt/FNwUZm8Odm28NiSQRrC13
aaiBOgZ1j+ommTMA+aMCTEbjCdE8Q+RDnKXbT2aJ5ls/C0EFrrm0TQ5lNkWzJ1mEyFeiXSjfOVg9
IrAE+p3vYs8a0M5lYxEZUoiZhTnPlcTpAHbmsQf/mDJoCGe+SmqyQwpl/A0AuEb3wQa3CUPgz6Hi
7B2Jb6rLvg1A98oZesa76np9hDBklMIhD+VdSDWa7LnhUApGquZVWdT3Gc1IRwPMW4YtZPcpUg6x
uqK8QkQ37NZ7GhMK7hAAMptK6WkBDtvZ2UtMCSWzp2NzadsxEJbGKAqCYR3fuL2Djf1D/9vkdth1
39KRRKDvJWqvw2yfeW6MATN0fv0qUWcGXzwah0VNSs5B5DTSbogi/ik3PdE3UrPzjshwQIcmyYg3
yYL6BvyxIoFtSmjdO4xD5EstF8EYvfpci1PtRGeFu+asyit5MlbjXpLZkDFLgK5OqfXGjs5Mk2ZV
RqpTKnj7WI9LIL82LyhRBc2mGpLiBIiX6tsPGVmj8G1t2AWxwhbELCjG20PYVcGNZWcGvkVOmx+z
pYTRyBXdGWgjC24T6TgLBY0y/SO1sJXjsZjJLOXOMFml7FIe6Q+mFuYNWIxWe4ao7tvO8oLKK1VY
qM1C5xUeZ4iu5bvbwjWZuvLKHEXXM2MJs0hTREuUwMtT1jIgspnlPol/1E7kkNeriRMg+QuCQ98G
nUOdEsO86yGTAABP7l/wjjOmsA3Dm9kM3q2Yyqu+V0YZK5Uk0gnXJpSMQ4e2Ff8fw4Gc077kjeNK
gPFTqp5lcLXW4ScUYnjtgm6s5WpY3K+3fkwqJao54l9Xc2dEmRsPpTggqhtYF/eKTsjP3KzQNC0d
/P93cUyJQp0t91mlZ34indqAMJzA/gB/gkemK1pinJvTHLOfutI5nCT2+oNGmhwCVWxCNAbXNDej
rn6msHZp4zneXYjWdaJEbWXhTMidBSytoEGHNBJrqoz12W0t97EjYq/Do43WK76c6cRrUZ9XYznm
r8D81ChMGImhlEzw/ZkMSCb2rkHf5q6d8vdlYHjO6HQeCPBjP2S03/eCjfycPc08r7Mv0g2Atebo
+mJkqlFo2tGxnxtlHnuHgysUHG4MN3RDIXQFaxlsb6vtbiqEGMTPU2K88TxXtncxmxMMkXGosM1Q
rXHKaKI57Mwxk5sDSBDEgE4cKHXXJM9Qmb1XUS+05zEytR1z1KiBEtjRJZQkWD5eRaBTiZfDGCC6
9Lnw3yzsD/CdIW4RXK9QHyfiR70IOGignJoTZGdvEjtgmrIJGEEl+H8nIjntmsbz4ZrECR7nE3+B
JV75fEMiAeSloGZSlRutE5BEkxxtbT2+lhloyIl3Z3RIIFBcFRfQuNj39L/UtfhmSJwzKEgtUbgT
e0DEP9HUvXl46K6KpdFz+o6HYpSn95yGMZFYzXCSyelqiPrciqQw7axmF3m2RE5jP9EIv6HwqPIU
mZzXAnpD0CFtMak8SxSFUCvhPxCRfM2Q8x8L1juUNG7aagdFkW0Yf9BZbZZWh5pNsaDrkmOVZhNo
QTFOUGJ817mLNk5/wVpKW4b6MMwmRVNdFa0KbKsndfO8iJJAQG8r15K0tmKoFl4eseX4CnNVtlri
F6V47rxR9JBqaJQovrFrFB0zBR7SacqtHS3xplJCqgcSpgPQf8zDRaBW/kx+vZCdVirFrOqebf/P
d4Rd5PK7a9Ge7gwaos/xV0S9lnh587h2uSAFjgjmzuYgMsqL6yEPR42ifiA28ewkMfsHs0SdiyGV
clRxtODyf6tgIPoYBRCTnNZjlL8PpKuGo0CTY2HJxrW2rsqzwPl6jFQ3jjg44jjQDNkgFJs4GhxF
+e1w2JjG9yF9RC+Mdh+jiIN4gRAaNEdSZIqhwq1M+Mpl/UQBYHr1s/DTjlVfpHfX+0JZciwiYcke
NEbozlQ2JsRJHdAOjyEDS3m/hgaOy8Q/G0z8p6HvXx8f0GRA2MV792yEJtRjjeH8p74J6PugA/kO
9g3jIMwb5akaEYeEHqAJWyvzyWd/IOuzcyAwh5HjHdbFOIAIwuFHsXMLrRfzTDk7oA5m6p7hvd2r
hab5hn+C8rQyF5GTn7zP9Xl3cFp5G6xqpWSe1srXlh1NW2e4z8D0MatNNUEE+wWPyzFZpbbCNLz0
Xh3N79fp6fxOk5b29KxCBmdi6mR1pGyMfRZdyoyQh0rGpJKr1Jeff/++H0afNcUuoa+feDJoCVIQ
705A8l4jeB56DVHf9HQ+5ZLGWTskyHiciew+sTXm1Bpet999iYIOJOPsLXyHLwQ5jCBEpQeAc3RB
+GkOC865io0VQF2gVITgm9QJ9AArTaliRtbHKnTl0lzYvUdBZqZ7GTz7w2Ox3s7yl6qbxaXzdOzS
T91JeRB/wbOGUMc0g3SZnYuHeCHpX0rzuKhgfgib/Qc21pL9d9WVAcDnvBDOT5IWxSdqXIVh7n+y
TxtBfay5JwEc8HH/1dVVADJoWgrNqrWr6e9Cu9xQJs1qpObOGUwpv9n1H5qJFKWHDZInh4ycMbox
nMRZiYUXehWDn5Z3RwtLC/KfxnkdlLVS86UKyQirpv8gVekMWsFtKZdQwcZEFjSGo3FJPPppfjHu
KoPd+5UOBsUF6yG559Sqf4qdBRfEFg1JTSTuqzs5oej2MvaSpEuVgcm33nhZHWfauCvRg5Q399sF
j3oFWYu3cYDZ+CbSf3I0AzrLkpyMrVUGqCdPyA4cgX7mX0YitaC7gJKVxtKhmv0fu26omj9vEuqF
2D22OLZrd7CDK0frpZDeYEhPcHRPuYFNGkxLAc8rHjEXVRbvLKJWvEoEYs2HoXMgvFHjYbaMUuQB
eFgVcMODvhRzF8X8gUMfQcprBaXcLadPTD2jTeSgJuy2C8vO3LeBLPpMMXGcwPj6Zh9v53UU5Ljs
cL6v0r8JkB9Qz2xyBc5SVBg9TmzGCaJcjAkumiJmXBf05UiTFaipJyJtSY43x8LopXdnTb6/0T6m
TocWi5sGm3wBHnCZdRoeHMSrRbCEED6DX6V8jqW2noRNJwMQ5buZ5J+yEyYl/xxPtpJ+xSuvQG0j
1igu0AeQcxF/Yyn9Iv9nzoRzzHDQE0wPmeXqy60wvzoZChHZOQynIwImoGIqtRggH56eryfdp5Hh
+xJAVyUJgEL9d3sQ/kDruk3IdsFCMd25oeOY+sg+PgAt2y3ZUYQP3a53Cctl4SabPE/7G3hIAsmi
tmApSYaeCBT1KXPNapO7o/gzlYtpeJ2JXjSDDwb1XLrzNWww14hRBeyjhyxmjhkBF48lIQIdGuNl
lWvG+V5QnYf8j7de9BbvbS/NQVyNARTZUjRxkexMuzDzh99nAFQyflrtILGAUGzdZdoVDlIftYJy
id6h0OOqOVsP8Z5ngV5qw3pHDa73GqXuhtO1tPGJq6a6JqMqaZkJQo3MyihW0DkSumr4+3UG0fVm
ydMZL0GWyLhpIp9zu3rxcdhX824Gz110pKQaFAw1ACwL+f5CcCvYqRpA1WceZtYAAkL9crNeCSIh
56XF4APe2QtAKPqilFhSsD+dmbBzCGOORpwzGvZx9e8bggmV86iOe113yFmKgO23+hbN+H+IJM9e
KiN0u+06ysexUcTIHuOPoQQ1s1T6nKiR2Cxw294W4L/fqgJ1z+tLQ6U2kAnbsKR8lvJkrWVnr56z
hrmFmr1pnIsKRjhLHCqII7Aaco7c7tTCJNpGytB6HeWPVJt7Yu4r+usSok+gIFkEKWBq1RthdO5J
AFcHD2aLdTrhflHAOzj8U0HLZ6sqBnM4IXKS5As6ebl/v+qARGQoMx98G63VMvNSNzvtZZMug1WD
H2H49YHK9YIZ+lr3QcCGtudyQswZiW8VYeey+EsoNI4gVKwLUoNMSISk2rF3CT8FWw18ojsQom16
gynX1n/vltoySGW030S2MTus3plM0WtCeICxj/rK/eAWIlLVdTtBqgnE4zOaBog3cJg/w06qYq1l
HHmBCcL3oI+9zH+WTWGrRzzyGoKiUczkCc6SJwQwPi8xEM4a/0X2tj8zrPb4xg9lEPH8Gk3VtYb8
m+rdSl3Pu+aUDbZudmJF0LQ7C9IPm7svDpFsdV3tr52qKEbOH8fGy/wwpJOGj+CjvAJ0l//9xkjb
HD5k2kbmSlyaUDp10EYu5QLKjuMR7evq0GYIIsEWa8pGBSYK0wux8RMUHmmCR2PMjwRSICzkseZO
ZyO4HPhEQpr0NI+WZRxJ5m8+C3FHxGaJproeC2gfWkoQTR2Kdqmd2jH91K7sQ/dz8oli3cS7jX69
1A3znRVT0mmm83gb2oEsuh6RXomsmKrfso+4hZJgaJEoqFxeBJUYdKaxrXGjEnxGM26xi69FM5aj
ca9S5CjH1uIgGKhBLoRRqUO3AB+gf7zJ6BgjgQeo05sa2majwOEfAgmErdLkKVA4VgF1OFNzw5hG
kPmbFz3f9zh9bOVzuOz8UL5IP+2BpDn8dIpLmMMEJmdfl0IbQNs7BDvAW+paORt+GoY/RDNvqyYJ
wIWPN0g0UiTQrxqjHoDRm2GdNKCydcKJeiTAou20JyIywSeuWndi5p/MgoqLIUNwBvWqPWYACXl1
u7ODCYgPr9lWBRp2N2pNHs8psN51NiIp8k8Nn/BFd6eRDk+zFJS4sjEZQFHEe9h940vP9CA7pVWt
pAPJ3WBLTQv8KMOm6HVTbKe//sGGIKvA/c7AsEh3dXbV5xaOnHTiCzNe2+AfEr2tFfhq/xaff9jH
jFK+5YGwy0EcEO5qOdSVSPu9DPNzUE7kq3r8elbxKP7+YeerJG3gmpWaTgSj01VcK2tQL6iIull9
h4suR7q9knFXdHQuPnsdO/ZSTEM9PU6FPdsfSGVPuT0w/bX4rrY6+5h+0GbUUcJKX9KJx1eoQUS7
FlzOupTgTq4hz/xuvASD1rEr/0PTy3Azgcj+UPkDDdIuZQV34fK9PrCdTZDDM08P/CWDMJXK8uoH
QrsqJM9IrdyAdSgv+Q5z2oA5A4lF6VYC50NRPCdrJT5mVEGxHVfR/Uy/Ul9UOepljFt5FtFWL4IM
fVq7FlOlYAKx820684QETnnXCRg+qpXspJBL83C8blk6Tu2jlu/8qua7njFLZXC0CVzSexnIdod7
K8139esV0tRpVP8Ju5hiFAsZkv3ShYjT6gLgnx4xb0wKx1S8LtA/RLAZCQ/jsJYoa8bLQFv01jR3
wKsUn/GISm7i4lgGnvcVR73j4VBkBPRZJCbHEl/Wa3HGPAh+tPGptrMxGNaFvDiIpEaYzAZXksGN
fxMItIOUd/U6tNPcQ9zutd8qzIP62eDMX3t1iVkVcRIwx3pI74zffEOP8sdg4vGW4SQhWhuxU+Dc
LUIb/6bjybpOT1NztQWcTO801HSXzupumWayrODUzNhRNFK0DAMAgP0PA6shnnz/akVQ82BLtp/n
ZtxclH/ihL42PPxZjdscD1m8EdVJXZhbs5xjVdZX8gLXDw4yWS7Tx2uPHeW36Y1N5nZhkH7HmUxh
hrd/TMEYVuAcYA4lWZ5VBP16XRBEmynASbwrItbKLDrdkqgPgO2W/UrVG9/2aCg+btCaTekFMWL6
0RILnJexS6RQAWsTziva2PFH64TF52H/dqtx5Gxv+jNdKMOSAR52av8gl6tZRli8t2BF377kMDD+
IP+1tLFKZlFS0acW3J5fWyZ0r754sp8Jnpp0DfoRLDilC12crEyT01Ax3vBQHklt16YT3VBa1Jse
aTJ1ZyfqAsRtwEs6zxDtLUanZPBg4qd2EDwzvHQP85AojF2HXlH+kM5JCc4L+jGwSN9A37gc3DtA
qIokUsop6FW0VNYzs5ravJwJIF980YtqHkrCByo7athxDCr3KXxNnTwlozPcE4yuqO5FnG2/C6Tw
EtX9McqJk274t/X1jWOkf4daa5VUYGczsWSaEG5NDifWrzogAsOBs2EtGDT01E/M2puz6vhotJb8
+TmPP6EXJPT0hmEeJpSAqVXkkl0BO2zQv+MJFv+ltA9UP+Nd7UVykWnUtsm++xmKUvOZUn3NAsAW
m4ity5yj3JlfzBlvUqo22EIAs5LBHScVg7d34XuX0NExi/n2Ob10uMhpc4N+gqsWvEObVmwjvsQ1
6fhv01cgaIZ/RU7/8pY4axFvOe5eN22mZSYFaxitykj7mAuNQZZusiwCE1BAu6rZ8SF4DkufCxiL
l25QxrXtcJqsgIkFz45x2bo1rL4xNgAaXypYyrSdtJhtlexGEUS892qnCnaHA6wODtQBj8mBqTdA
amsJcSizN3GSutiSTgWRVVfHcAi6NW67H/+1PQDLAmJq6hLjCBqEp0UvbzFHw9KFTbUoJybDpABs
b86sWohoOcw9mNdgyoIndnztezBC8L/C4lqtaWyhp17dreob8xv28EFOaq4ICi+7Vpd7e6Yszfus
9KBL2wmWrQyC24wBLEAX2sytA/N/tZtXeCIkboSIyDbWnNWKBaR+ad0zXTrX3sh1vtZmN52xxy9e
hr/3XyRXS2KKFSUDD9g3VtJwcT8TXut9+yLJauS3tmBLAbzGWNGMt7l8jZAAT9n+E6HgZ6sYtyU8
zGcoLArcZjOF/2B2YkKMrr1EHTgo+tRbxGD38aXeH8dftR8p+sg1KWtr/zqEoW7wXUFgwxHS37vN
yWILidkkYQZiMbDu5/GSNljWiJDHzL7nNCLras5mPPmniSHIVLLzWPIMAcuUJRFvJJASjo8MphBe
UQx5S9k4oGTgNjT8SRaeM4VffQQOK72VgODGQPub9jkDnsNcs+NptMJpV7ii9OJfEXXPO2evu0Z+
okL7pGcp4g9f5E7s4uOjbFJfS6PBcTQFzmWosZGcco2yikatbU43rHtFWh4dgvvAEVNILyFDz5/B
s3ZOJ/b5QrmR/LmUsSv1x3UIL/5p20PNIQd/GfdW3m7DyrE+9F6KgAN0JWk4Ih1DrWBM9ZiiuyV+
CW39SmYEsmr10NJxGLTxo/yOpFVAsVDE5w+fmzhLrJEt7BmupqhRpuJNTpwalh4dIDBS4sttGUz9
Jn/q6RMf3B3PqatXKvzewrIkJvyj+STslFH5LlbIaWfPHo4kFyA8NfyOO/QFyooI/HCD1edHvBg9
pGYy57CPJcYTqWct2eoHOgfa0OER6N5fDO+l5CAQEgf5eONO/2wwbbe4dUR3r4ujJPOFkIrLG77W
D3QBtSOt7drNISD2SR8T+2rHrl/dowANTGStWDeEh+1C0xGW+7gvDt0MEhKEUrXWXQTG56EcaeJw
pQ2QnClz+S+YeimphJFZwH0qMN4Nx0jjQQpVFi4VxKGswQ8bLUk2PdXxzrfDUEmyNoXiB30xt/Wn
eUxwvGigUM9s5IYG6ZITcwXKrhV7nb+BVH82r1Z9LEZUHMqaeYAwAWFV/+cbP+ZzH2NBfxVFcx3B
ywm+iHTMr4hGzrO7z2EW8b2OLocl465EPVR46qFLbCB3fchFfr3wqGRZjyFf9Isc+kwBFlIJKlSj
OVxc+jqC7E/ysqhFBYM1rnw/qrt/ujkaChfQGd/PhvHoqF5y3KSIzgqgsPhXdtnw1jPXBWII5tM7
D29RNrIJ0bHVQyIwjOHRALBlgYSKT9hpWR9HnvZXhzHjxZJap76rB5iG9upOde1MZ6H5DabbGpay
0JCVcvLR2l+ISoPmj2sobUp25r1sesCIsKEnfC07HnFbpsJNIUARHUU5eHVgSnRJLX3xUDS1+DOq
r+oC9vg+IOPIg1ndKbxLO+442R/OKfod5S6w1q1qVPgWJXOOQW7GbwG5AjcSbRdByY5lOmi4ps3j
Kfud/oyrnx4i7WGQLSZGMunJiwMV+q8xnTxDU+qQUfWwz9xOziBScaQfXrwWPe6jx5xLFJx/PO7v
6LXPEIITe855qmwUEIUaf3XmYyyPmxxsfX2Dxbavnm+IrE4jDqsaTjp4krUM+tJDHQ4QrIX8Y+Vf
ldtb3z5Hsj+PkyCY/ANhHNpLT404Cc/kvKKz0tx0BHnNL7hu1eaU8fltCZYjHLWzu1cSktY78RF+
qQ0UEzHq8W+DfZml6ZSPXR3ZNmn4UIKsXQMAXtc99sYT0ft97LltgeC6ylMq90YprNpNcigv4wZb
NHUiLLX9k5s2XBlltTKGRAQAIAzCuecA2KQmhCvy474gwxdzJvwZLXfe3RhqVxzEBhFNj51zOubp
6HQmpVn46+nqqPIWymSKXnV5giT8AZUIxzvHkTzS2m83aC73pjl0NG8eMrYWerVkB4v5mbNhqOhB
KJ+5aHALE2EGehV0snPkpBISk3GGHXqC+6PcVWFZIPVJfyVetJ32bTqJWooHYoDFDWibX+90bQtU
gqpxT+sCR+awWg/cOpRCUF5PCiZg1Jg3urxJPMeNgP9PJ+EO+3nC6QJrxDwSbU5+/zRjJ2KrhP41
I6uRFo3BFz+2L9i43w1te6fCs2keqLcIUqB/c8KtRw7/Xd0+unp7rNJkSKwvxUhkD7K21Q1HqmpF
3HgBwSg0LaIhy3aL5btI5hCFNTG4vc/oyr9PNTno/fBEOCEnovk6mVHrKEd9Q/Pd5xutzhKsdk1y
otnEeFQPwUhgwssKe8Sr2d86wGgNQg6yLwIVQSlFPdb4InhwAk8AVn1bg0HuhrxqvG2mL81w1Css
iyFDw7CwNyFH/n4vlsNCMRns7qoa0ndj8Ev/5I9pGk9nQ514VwVwsof+3hkSFuiyyRnskMk7/yvK
xG7vSCFBMOtk1RAx83QdIe2jKESmkgVADe5eblsVqxN7z+Z2c2pnuPK4tm/WwFymL8a7h3e/IK8i
Gd2pG3FJLNHAlVkTGLLz0QZyvJ4LqM4CYU9qfuczXxpr6KAOtrGj5K+zU8ffg8Fzks0e7U5wO30e
BV1ZSUWi1hxEtgty0qckDpNs98ViyTERrqIhbK1RulKi2OKaW8ykgcZ0wFcl1mbdEZJB+3GRaX5q
wdfIxSfDe7xno/QSiAq8Fvy8rykJy8u39ksGa+UzWhoimU/G4i4JWzztVkaHD8n0zIP0itV236f6
v/kCzHsS8B05ZJB1K6aC1wgIled/uMTWMv8UM9V9iQ/CkiUnQSm6edbsj8Ka/8xBTPY5TVsQVO9b
G0lWQAYiPpZe0w0c1cuwKJc8fEZUOD55VYmU3pfxOSnVHvCQkWlY/LrATcaNNyNHXvNo5fwujsGU
/+PmO9Gtgr02x2yhsR2eEbjY7QjG3a0hEnUvJL9g0h5BkzbbFJNeKec5Bm9ykm2LaFW7RRx/vDgH
q9WVnCObMJ71JPz2yHgkliEDLiZimWsZte5XJMYaPBIh9x4Z0m8laMVVADnezs4Fnw4h5A+fe8pf
4KEje2j+kc2D4ReTaxo5+ex2rwEpE5CG155YX+25jKoL/gmI7Vruyk+tV7uJpOU1b0AD0mjgOmSz
O1Coyrl6vmwboLcvFWvaeYHF63FLXOSIS6dhcD9/5Fb1f/85HRmtmr07SipYeV1xATsec40pGrMI
R8TjsKARGpHJluweLjeXSbxS2WzLLeR/RV9w2jVJdsCD8O9GKUi2Dm+Wkl6hUm/8ecG7oqs1hk4C
uxaYZC725Bbbwghcj/bfboVRdDMeWxXTLjQ2+zOfboXc+ATJ6qwfOKimm2Z/zb2b/JVzhw2sqdqh
/vpQFafb/wGsDRc1Sw6oB4LTud2mKIaDtG8/T+rpbxgDHlfD2EPq1g1IKAsPp/BsXPcHdDutAMKX
Uc0czn6C+69M1N6AP5mhmtdDhIw0LP8/3eiXiYPTsnLodqEggjPEdNHK23jSR2BDTSkPXgPVnRRw
9jQFBv0W/QUt0UXi4pOn1nmrnr/ev0tUA+QYAgL3yDuyx4zpaY+WJDcJNV3RCR0m0iKjq+rCHsIU
+rKBdfqa5N75Rk1DFIo0HbaJE0CcgyIHnSJnApiQa7UM416RQLJzRrjmoRLOHVcas5uHOiYuT5/6
zLgyZgTwpTYYbcZKdiVDKwhrYTFluk2DbWrjAKYw1jsFJ/gPsoOTYIm15jy141AGXMo6kmn7PIdv
HVkzMmX0Hv8vJru6fyDzy8V0gde388V1OJbthY+80qxL4jaZv6SwGiKyrbljJPwn/cTj6Y9qhUES
KcA9+yNYhbQoAVP3P3HjNYSUFvF2Akh0GNcumeEUWxN9YORQNmNjpRW5erIjr8F/yt2/6K4v5PyY
VqFT8WD7RNWM3aH0wRXjs170F4iyXe0M3+lc70xW+8sHgi/Y6jywYZZ4H6sfBivUQU4YI5Arzq6I
hTDmj9ZJDhE/HNT3VG4kcKpZEg/cf5JbZ43aNghBJlTzYKcRdu0+ORKd+0Whp/Xbhyxb8Mgkf0es
YLpvwxsLCHowCvbq0h3/xnUAeV1+sOqS0vekLOaj2J+8kjegyTwuG6tf7TA7n3X6cgHOC9+tWWmd
LqEWG54ZzcyHsgyZuF0Ek4i4moqX8P1ZwIq2FNCVS2kVNifvQzynmu6rwGAueTx3NpIZDcb8rJ2o
gqTsKI4YgY5WKSXO/ArxorAkGgC4fPAxm3qjcziFYLYULwUO6pPhsBrVLJVk12AwlBUK86LqGFsg
8QnMzLfqCf2G/B8mdcuyWXmxxcTRnwwQ1u9LROOgGiXQYrBCCx1M5w018tmm4c6t8cx8GvZ4+dq0
x4dy3hqIZkvFtO4WlOw+N03xaj6Itd940PBV2fVQ3UM2NQrV/7Udoas16a3O8ldG9O80cNl1/tnX
iBmLq6En1UObIIrGW2eUlJElB3NXT0jBQxffl2lyhNqnBYl6gK84Yg9JOOKBlTjHO3ePQPXvJyZ+
2iZatyHKNK/Cxs567NI6IvKQoGXSkh9KRDGTwPYl65SzdeHM9aVvl8HQVzo6dwNB3/CGU3IfnFqC
tttTjY7ufm8JHWryUxIV0fAMv/uLY/ETNRI71QWT5FUiUELP+n+9+j7rZ8ZRMbVyNnboJc1f9r0e
5MyCR1H54vJwVgpN3pMdOGYYQMnBJLzwN4LACjGcAZseBcTGGiU37p2tRWPdhYtRhDTjTJvZADb9
IP1DlBzwIGnvsGcSKKnL5xr15Na747Uf05N/PRmS9ZuuU0AVFLtegSxyZtE3LtXs3b2xYIvudZQp
ueqPFJ/YL03nKEy3ux394zDXBDnAqLR+oZwUdtIcqkXymZWiRnyN7OQ1LpJIfPVUhG0dghR3UT73
Yt/Xjxmm1CpKIONdNf+NZTPloCxR6fzNM7HYxbpnZsHzHK+BDRjO1Z5bGp8gNhDERsAyetFyO4fG
a3Q+rHXavtKKV/EawsVhYC38Jq/1iP+5DmFT4revJRkoW6oc0W4TKl9/xS8mcBv9Z7SxSqR8rgGa
k7nFK1c3z4t0UY8xDml5KHz4yTjTDXzd6uJ9yAt3xUUBZk84H4d29MdN4GXttaoUWTG7X4mQcs3Y
w8C2xneI19HswW5PXurEaCfuFZvaS9/NhRWbND0LVSugYUT0n98gWQG7jxQ6+obuDf1HmWLKqbZR
N0GpR0UDIYJxPJtYhRcwsr8d0D408UsEQTU+w0Ups84JuUbl2DB3paKpnVaNIj+b/O/CqhaBD876
qa8YX7DckoiIyO/iIlN0oRN81S/36qysTcUfKG7RwOi14fAnOq8IppL32nXIvEG7YpYbN2/hpIsP
CV+4bjhby+WW7vJuKgDZDQPmJC+zgeB9qiKmswOuTVKMfpwS7z72EknxcdYfGo7gDiiDRJwSpHtM
a2uOLVBIfW3NPlFRHBYhty/jSVR2FFw8/z7lSRty6cHmmg82F1uZS+hIXd8nFrUWvpJ/CfVRZoF0
A5eRQVVNZfAjd1rRi0xU62Fu+zwoKurWv+QX5b9DJBSPWE+r00dZC3jXEKc2bHqsv5+VluZGWhVo
7t0MHCMlsu2chfe9ir8oizWYxEHs46MglC8veNO5goRiTOyD7e5+Lzxxa7a72ZrBuTLD8xTEOvdC
Xa+BWiKNvbvTfTJoGppdUo6yIOhmpw7WvOcNdZQt0CL/Kb53/AxMq1J8UGNE22Uj+vYvrFy5YHIB
3o6kOFS0MssJ/PzvfoUGBluo+6adCdJr9S2LEgLvi2OGDzbcQDrFfgWlqYzly8RSawrsMR7JU3Ls
uksUm+mRbZOAFB5vqKbEIqF2tFIaFtlDurslXG6i3IEqTFjIKhl9OgIGH4O55u+rfsYz9V4Mwocj
EJUaDNDVmdFTITfP7Xx8nAbPMW+VuUHyK70HhqBL2UIyfntpVYJ6BxKakNOjIttLNoBuYhCleC+x
1tVcxxV0sMv1hufx2JqzvDP80n5Fclgw+IHKSZxrHZHF9xl9h3sHZCRICn6Azm3VkBuYalvevDoF
wlRejKi/fMwvwVJPmy64M+KvoIMU9OxI3Sax/OrOE8pvp6cJfp+xZ5VDtfcavJ7+cwOy1vboxIVN
9DNgLRGLlvSbFUEakPEidgPAT8/YbQQX99LvClDYZQyUvniL2D7Z8piRrkf7cAre5860/gIo7FTX
6CpikDulYEOy9q0TI+Swz+Muph5whXQoZbayrBeMvh98C74oy2EjXUbVuKcRyEn8a09PSkx+/1/D
D2ZgZR7eS00DBB8A6kmw9knPkp5KBTp74vXpozaLQKZsDM5GtnUn8XP52De4vf2vblSUTEEt3bjV
oMslsFcadkwF/EHEbmwUDs0WNBtKyVnqe+XOv5ID7jBZ5Q/5saBlHBtKJGOctkjzNJOAAPgfYRcz
phvrDReX6E/jB3DCUmHQAyThDp0Kl5RnShYsc0unEiIs+jr9D3UCgvA9quD6fDAaxPekyr1yRO2h
t3PMgIY9mO+3NZmA9iLe4IqKVh1yzIzG7WlUah4C7VJvQU2hk+fjhUjaN2SjosFcDZmHf12xq5IU
K1nI4yIyhUhxpxodnFxsGVcLE63vSm4QBKTZbFTEUWnVGVgOueuivaLvpJ/yT9wu66PoCb9sDtBP
B+/oHkgiKqwYdo8MlwY7MGZIjfRP9W7oQc59fC8D33iMlP22Zo8e3B/IxVljH0OkhQQIfDF8qVoQ
nCe7SW/2tMmO2qSCer1q7Wl1w8sM8Zdd4D309FoaJV6N/4CzUQVWPfHfkTNA0jmTJYBlcMBliusf
ydXO+rUv1vTySX4LiIfubWigVe02GIxqE/N6n6yDE0ifZ7zrmydI89rjTW0z+WXKaSTUFIsOHgzh
nDYS29dyjjY3MIQmuKvazGc86MBkO9T+0gzh2zLHJm+8MExL5hWDgWUltmOCYusjyWzDCg9x/asq
qpg3W2gHfT8m+deCyb7ZaQONmP/Ok6rRFcaTw37lAVVIaWc6ubwpBg26ThIp7JkJWfKBXtRN5zkH
hMZA+8wvsK1bzxgMJl/VB0N088BLGqgSd5R+iJCiBMp+eKqaoFKgcPwSG+JCZZ95rehQVyF/QRub
J3VVvr1irUjDvIFbDaVpwBTLbiF21GV1JTPETL5dewTO0yJjNhfjzTKw9xyRFNT0HhwMcO9ZhlLd
gJnOQ+ajoBWmAr3QJYKTjjNHoaJtpTGgdnkxG/Yo4eSMUh/gIfs5nUuRkHc2QjuUZFecjpB4PvmR
svGmJiAu2azSApAo1OH9go+pBEhSj1EBwYLnEaZLYT70X+uxnMkuCayAacGJfPpPDAKrcPBDPxrF
jlGjonk8pg5YbRyITm3hpqyVtRKNqNzlD7RE4wi7Lk17cVm3DTHlQx9V7vm3VMVLLxihyhFwWRMR
W7iy+gL1b2E7oQOlEZhOdmvRyVzcuajgC4nM/f0dskaVCY6RKYo3oUXArq8pD7+XX1H+4mpc8apE
8VDoWGvlvq52KoIhBSFqYxY8C7juppAsNpoZdJkMfy/CrQj74zLZdvgjvHHrFD77FK9iqSmedkI5
G4ynaeEGc/VJY4LaW3y0BWXHfjHAYRrbYkUJYn998Ed52sJXXeJEPgR1FO+1jR6/ZsWWrnUlsOvR
p4h5SGnCjz+QMs3jMHr+otFk86bPuxDy6G89oMaFti/sFKx0xVm8ah71AM1PJqlXrPTSRZ/sjo7G
At/MuICdFrj0cJyzekDg0av+hYHw4LpJFCANDAfXJr4nkpJgwUPB0CscKEYkH1WKjImCkOYGRspT
wP0elpzAr7VFyz0l20hKafAIQ/LOvEefyq1zVa8xa4nQs5j/ubfFLeqfX+fIOpALk9pXTgHfzorV
tbYqa2JPRi9dSrudAwHSEUNOq+gCCTYR4fhFqibyCtIsxI4YDU2n9cg2oCbZ4km1eomqpwy1xdwF
AWMs7yx1zo0jRXvjRUX/M46QlG7ZJCROXKZ2/CPN3wct50d8zSE3B1so6bxKV5IVKGXVkcLZNyhT
BjUlcMiAIiwoJ1pY8ynsciZvYBMeXwvRiRw11B110bqJCYqhh7Phx63at7lz2pOWxsPiQrIVbbu9
Cn7jEgeFkQGzuFVQuJsh0raFCxC2CW48A6g3GMsW99/NWKiNZOsSIH3M0EJqXYBp0ogA3E5jHCOb
0CKA+llLoa0L2fFkWimZpwrg6TphfyCyFRw9U3UtP1V3/KkL/OUmmzefuuG1T0Vf92EXT42rlWx3
1IWxoA/TJVzYI2Bsb8RvoRoJgoLBq9oIv5sRu6r91/Q61oCVRHAcuTW9BCCDUxyMgNRlcBRDWJkG
BFVDTq1mplfejQv/S/fWtBiyN9ahvCf6jjOFHHlQ7BfeqVgaMH1OjF3zVUU1iGLcgb70xKf9JEN6
pT46sRmZmHovXp0DUTrDFKQ/JMYuIbHRrbvj8FLVh7qu22siEgWPxjvjfkcOnu/Yoa/pUsB0eyCU
U529b24/HpyWd/ZPsCpKIGm+D+AnVo0QNYoap1dhoeNd4QC3psuAD4hbcTOZil+uU02c/2T8VFpZ
t0N9W7RNqrI2l6jxz+og3t05CC33S/omhXRmuSRYv7OGmf0q/2qaNr7zCI+XIdMwNjHhasFkL8VX
OfSZ84X+5QaaxgG6dYAzzJ7WxfcO3Q+4JDjwAJ4ikG55f3SRWOdOxHpG1ODNIA/HNOI1lVqi/3b6
Onm+cgopvRVKVpOOupQmORi636VYJ5qkHh89OX5/qDrUk1manWH9cNw8PcA+94NMXn6bedJTBBuw
91eU/Rg4mAaMzIEJwqhY5oP+wbx4Bs9WGzzkZOmbdZFVPmyNz7o8ceCLHv/p+TJdyKzLKFwBCGMP
LOzXjf33lnXCRbJVYlCsceww+y2paX9iX4M2A10sb3Y7C5kOKdCsja6/PkoejqFDWt2IkE7V5jN7
u1jr68djwCsaJ/vFEhw40Jtcr7Voc+WseRJkC2HzFuPEjOhf4xbpfN3riE/tc6wddoy+ox9SRyaf
GZ/rM79g7HcJeffZf2ifkeCQu5iwaJMTuNvTeFlM7rKvJydc8LMI2EF38WOWQRzHxeX09iTO0UKz
czew4jHat23CPALEOrAHFtxGVhUweZZMgtFY4LZQD/AAA219Adgith1OP7GKno1fMmF50sx7A2lK
LQMqQIENQ9mg9o87pcHrLcqBbNGnSDsDEjPjWtmaZta8a/z/xOFK2yVnKQ9yHhaWojmLXwwFvRCt
xG1oZBNjKyo5GT+54Z4QgYu4kV0rfl7uj37eF7C0mk7tpvsjJGAKGoJ5jFITI24AqKtpw59TP+cq
powL2dypVTX3baZNBRVzjcmPZcYWnUy/QQvLMwo0WNrZF/zBT4ClqB0Wj79Zey5G4xS2lfvO9scC
nkr2sFNSmd54bIERH6iMxqye1OeUvJsMzmKZaLDXy5Yplhzw8P/7U4neXWpS+WvxtWVL1djgaUt+
qosj6I+iqzIJeNOD41VC26UQ3QwW6oswYhSeSjMEoG5QaHPSUbBAHTA6P0pE+eEwYJDnXAP1qiRl
ik/VXdhwbVcWqK/5gWiwCNwY+Kpt19RHCm9Wb9lTaU/lpaFzmdlF2ZO9DB3CSruTop7PvorP1dGN
fpa98htyZPBbbUjOj6pfo+Q6kQHp8Zr/BP9Yinj0E5t6DdOraK9MR2b3fDdR+YVs7YbJ9OerP523
rxs3bkLbLaTiAsGWa7m7i/T4A20mdgIJqtbi8lUEjg5bOmGpqy3KdklH/Jq7137C8bB0cMkruAXr
/TFRWwUOHbcYMTYqw9B1beUTmfrrXUwFwKXn90x7hWCo8Xx55eG+v60nSruqx6qv/ojo0ENkjVvn
yfUVroyARPGmuRiZh/cdKVnCqATVEVLARS3G3VbKH05FgBF6aga4puopq2sDwP4Fda33puWpjYUb
NBVIPGTgNtHkrnfkJK1tJrSjsusWGt3pKowFmH36X/5HaIfzhb+OyJUSMgsc9YOvYpTAFIAaB1KY
ATABLnGHoFryr+FNstkODErpIxCLPYSCmbu1LsYsMgm2MYtpSDC2/dvR+CNdb4i+VmIB6a2G4lJE
wL9fDjF8vJJaanIu0kX59f3DT4QZuO5dw1bU20TA1lo8GZckwnJ8GKtWtOQJ1lOxQH54Daatempm
SsqbHoNXzBcMma/5VpAEg75eYVrsjPNK+0Co/OLu1XdAC4pL7kyldPONhnp51E+yhWlWZYQnOzKi
QPm8QuObFwuQCi3IcrBk8QxTUuAddzr/A+BnKOGyGV6wFj1U75R4Ob2c73kEDIirzyXrIUBvj8mw
X+zE5QZJEwEhDqYmDiGoO64FIJDSSiMJcDd89f/4RKUUznMKEL+dKnXw6C1NlDmXYALIMMcl5u4J
ShtNqotpw8+WAyETuX/ArcQ4quvVXaydPrtx5Ix3VYDDqRh7IThgFSUxb3sOq7kNiDHTvURG94Rq
u46fxriJKhCHtBAzJeu6dn3hkGvqegORxGQFMgK2pI13HpG/wKyoAXPiFm1mpNDThQzNg7cSLAWo
kpgL+zroeVqHE/VbU5DL0mI9coCP/jcGEs5/fxUtrGCAx3UdaDiliUhqt9Hba7i2W75iTxuyZlCb
L03Vvsa8abExAlSXNqM1Y/WIoovVRmf03AFHg4oPRaOGqio1fUeMQBKGVSc+dDQXrDCAWynnfpYs
vxQqbBzGRkkalpMHllrIN8tMSdPOJ0UcJApC4BXHsn2Piv9gyXJJMpes0S9hN8pG3jOcuwC6CO6W
bu/lw/+nWeg7oCY4venqfP8hZyv6FvlYbu/W7CxhLw0A0VRDmcLhYOXnp6Pgx1VZrjPzOn16W3PM
9g9ga448B+Z3M2gmJP9Ndq+Vtx+sdmSwnKEviiudvgbnd0hiO7YZrOfc3SC/Z3oh6/BkBDjZlMYQ
Gcwo2nIFDuE7npmSb25Wi4edEOvEdSgEdYMZ9mQDaMcXFGe7fN94+zYGZ4kOHQNsYDTn0LWvBgcd
saunJmk8YljZIqZrNaapr53a9LgZVZLYhmLoaL4QJJUWqr1JMgG7vv6GR/ggJRaO0jc7X0I1E4Ux
Sirqjer+dXmr8x/KbOlEijjH5TCT1la/9IVnIXdaBd8zjL4FvA1mNDbdf7UrgiYKry6F+ipEXfLn
5q7tTAnpQiyIWm6UYM+BrELOy6QOZvqtLpC2ri2uQfHRAe04cx+cb6djs7Cys5yr9m5JfXmOjPwz
0s6+bgmz4oPDrMrmOoX1VQMx7ZROqmrT5rhd8dm+hLPevlIblZP85vqcHGFuNL2D7yHPd4FWHJvo
bo1ALQSPJWiRw90rxeaOjQ64CIVNGpeSbEnS3iCkun2LsuMXcOguP361y6Ut84jzeBZtEtI7iMXR
iaBR/zMcCUGD+GEM8H48npC19cS+oP91k0ZpwzqVkISkMdDfYgnrnvZPFzqSZtk8Us3aLUWKLTtx
9IewswXbXNqwL6jrRE/m4EHFYIAa+lSAARxUFGiIQjVO636+j9hgAka3JSta0p5Wzal2XHunkGN2
0kZZM3+HFxuEfA3z3ZqQtM7EOSBFR2XXw7srPFsLASFLI+7bgeh8xtmyhNPOO5sVQ9su9s9IZAap
JraJVBeyciB9ntba3UAItWnCMQEvhfHRrRIBJTFdwgBagbipTjmLDi21+skSqmcCJt9NbFUAUHXS
v+r6lT1HLJgXtqN/UCYwin/qV5QVqvFeaFRcubipVXOp0qzNRWkIoZ8f7GsIidYfLo8G+KwiiiRD
pCMuuaQtZdG1b+HabBhGoMt5yUIkurUselVqHf4wXEZuxiAkY01s4YUXLKv56TntLqkPJfcPT5o1
o0KcA5VC4gxtZczdoL1947cIEsvINeHMwN4VttXscobF/ZU/Hdjubsl8t0kzD7nj9+k3/6+L0FeT
2qxg/bWru11ivJNzY5R9GZ8Jn/RvT3KAuqxdRMuSdAqrn99VJAvLAxSlej6P+gijkJSo/e2NJXGv
nIK+D/ziZswyhSIN7107k2GuPj7hrNjj65PNBzKcfh6Obj34Wz+anszU4PGR1gKl9NNtJ2th/6w+
m16id0sxDYIbQ3/5Gw3Tgg3VGHozqgMBFw3M3dyV+GpsYCPsDho4i/8947spidvhuQvku6FgQzyJ
eQtyW9ac2E5vvReGirN4MA3S0qxQqhpr/krs7RUXEaggdsDlP/TFClgzy27jivpL07xzexK0ksU+
3lkk58wwyBTLfjACE17XV6tTzK4sVCL4yS96RNEcNI6wM9o8Ao4wWlT+VEzU1KQ8gp91s+6jcDSY
ZdSFVL2SK5IOgB/RRW/fKmIGhWuQGASBTV8Cvnakx4e1BhxK6/L6CxM3bBgKHAP/9LlNI1aIms/5
e6S7kbdFhj1zHU4t0Gzr0Z1qlogD9M97UNUSTohvXiqm8KXRABx93SXmKZV8z7+mRdMdi0xGmtvX
p2uawWAWrhllbah4j1VUs4UpMfAI6z8HJ0KUkQH5/cBj+yhWiSyd9VFrxG+1BYlqErSSWQG/1Spg
QZCMks7kqm8xOdlKFOVl3K0VQAvzeXgdebYVKOEJONW5OcnTbbfhVFDTQGIy9GVYO4ts5ib4MZUe
R0+Da66t9fTC7uSJZ1tCcnVB94rEQlvJAgZUIQ//92uVu6EeYbAWPQ+vMq47a6Rx8hUf7kH66rnb
tY2builhRUFnXtrlZXLCxdH0hJzYJFmtgNkDo5HjXIfBBLqYkq5WYMHX8x8Va6zFVCIwcVy8znZ0
+ecu+2wP9VnNtTT3EK6RTkWBjiFiS2cT5YkbhckE0ccOoauxX2RDNAZoWmyAnp4uhTc2gjBSLj0R
l0DKOXasPdMIePny0vmmGqZ+vklibBf9MSY3y1R+mKJ9TQ6HgbuqTW1wHKByVz55qZqQyZP/MnMb
jJCFmgcvGbQP9dkLfklHiOd2No4ibUE0m0+vSS0WmuUFUxeDPnqZYI5H9hWlbYrdFOZhWtEKJlxG
FXXLnh1L/pCZS6HTrJxBIyf0Ya7TKEqW1HgsHBRA7vcco7QPX22nvBUvS2DG5B60Ptr6yU0I9xoZ
wT6+RkKVmhGv/ffa5aY8ORMWVvGLml0LVPkc01oqxI8w+QaVFFKFe/mcy/NGErkt6fT0VFz8aa5y
3fpa435co4hh4g/lbq+P7uPLAMS549GQEsbhwhjBVQN8KncJYeHRq2wD7cDz3yX2zB7Z6fWZOlGz
enAH1/jahq14DaaCjKDiczmTZBUrtDjKDzNeDUoP2CXqYAl5/SGlAfAUUloTL22ov4WXNnYshjqd
72/OkNMlERsZMQdyCzIegOekS6CSvqDiw1ZauaK9Mym4oDMCHgHaJb6k9Z8S5aoK2ztEDt6wn248
MQ/RpWr+Ib5M5w/DTxmWEcCu/aJei8niV2PNrcEQaBQ34I/vJtY/nDbcTFmrSeAg3MnPkcIMamfT
GDyT+E/EMffE7KcpNlGbWjyISZLClIn91bzqgmHtQBo1Zvh96Nkt0lH7pBzvqe/+Zwwcsami6tZS
Plsu/I4V77BvopfBiJRtO/UGUuNXtlQayuA8HfsvNdCMbBjDTDz+TYaUIIncYmsDA6a8jQAIyhrw
iU7RitYNrycbfdPBpDWxcBkVsPo7+CSa9EKT7fYbTE+tR6j/1MlssPJIfqCPDvY3xPZp8GZCJS4v
xhKW83Z/g/17ljZVTOj9YpNgXyWQhPPHIeCE4vYRTnWfgGaLCQQN0Pxc0hUh1DSma3nCI5SyIaUF
OtgyoyAc2jsm6etqtaTd7+B3h5Tv5f80KrTyUDp5PYzsNgWfS9RIYTEG4r4sKYXsoFNfADqXDrOr
fJrXE1saQSKP+nwRXnx/FTSqfYodI+ebtrA3/sLxG5UlZ8NqtawN8RAnLEl8qquhsTO0IPdQkA9x
f+tOZ1zoGZzEfWl8IIq6xUey22oB69xATyVAziLWxd7om7xRlymT6bBW3+GjmMMtg8U1/k+atd8n
GF4gFwBiYXT0HtgqJLjQNjrhfuka/IFj42Shq5QSvgtNHUcR/M0XGjOJscUtEsHiIqPBv+aflcoR
t8IEVDOuJrENe9sAvqfAXNkKoD5PkB6MVDyZOod6LlfJ34/ITZ3FSZrRgjV35gnYKVN+0xs7Lssn
LaRQm+JT6kTaL50maSMTvKvh0G/UNn4RYe6NCO4RuN7SUU/yO58rvd5RWTBhrYq/Dm95CkmvNCEf
N50Lf/NuCFtG1Z5x7gPrLZGFuC3Wv+BClj49QTIeAuQSDBqi1vzYSkBkn62rwRmhNlARLAi0TTD+
UPYL0OYHwOFuNTt3XTxW+GCGabza8XMBebejTd73LCLvZQ1oKAQHKJewfXWjAv07jZblX+cyHMPE
/Ds7CwZn6jh/zrmTgus5dYm+HIqcMc19e075RtACgLJKIa9OESjULned3rZBU/6+1pp8tfB56OWn
NeZEJldo3DgQcFTmvVwC84hSDj0p0MKR7RmUAVD88rDcQC5+RpOeJS8dSlpNcYtr16Fb2ovUY+sw
QxPqWNOzYcQ79IC3GAYeDSLCn589BUCf3Ew490Szxm5zmn0wQQb3BBTQqTJz1T78U5HwdJsIYVXu
Z/01kRoRmwO42+itTKk0dmB0D9cOEmPl1vk8k5VMZMkzd61/ROt49LqAtfRbrVy4ahW6L1IHDrHr
rf2irJlDQWrMbJiAENC/eiosQxdStqG+1e+jw2n1gvferi3jKw9VxnnFms+epeYSJU3ah+/JIy4d
883p5rSguK6RvwgJnzHxqSt2Ar/Rz6W5WyH7M41wQoUm7UnTi+71n9Gqt+/DDw3w+yBCamrfbd8t
lyO5v+x7sNno1HAdTsEMQmv7JKMMDVhlJCsxzPaf/ylNrXmBJI3anp1IfAdV7ijomXsoUiDJpiEk
UMzG57arokt4UbzAessOVJFvgIl3tGrx9uKeuAOWQeN7BSLF1HnHSjAqwRVDl6h06nAcKSZyNQcC
uilgapaEWTAOyNCxUnTNjFUwstjxZXBlkc07pVvN07qQkwAA/ra1Q6IHqDLP9M+mMMMlRgkkiCp3
kfx9hA29HXRZ7p0OrEaEKVITvB1KyGDaGQYA1vc4ZzNjlygRi01XLAKviZX3W4pjQLkjmAlnZnLC
EVObKVSVOkKxDsjRXUWj16Yp1JhNc/zmNN/mAPcWQOiVQkAZ8leO/XgA70F4WoR35ds8wvZq9PHs
D6avmwqFJKe/sukSh6wfuHBA5k9XfcneUkFjxSXo4wQOmVs8+zlVpeqIzDeR0SRb/eANSkgW24oi
vdJxMjykzstI4JTEzKC7hcLlGkNeiiRCPZVVk3s4fOBy8ooeFQhuhxWxL+8/wqM9ts2lg1/3lphG
U5kFPh2PCeH66fxbrJwEdFxGWSKfC2+cuVL5XiVVbqkVWwoFD6DOvWpDMOcplDQXiTjMudGSxIMy
ZA3Vw0F9ZN0unVCehEciMKCyFrSYjxPxPB54QKB+FuvXlKfdUoyPg0ualR0S0pd7h8b8LhCPufOB
hff0ZYo+riEejF0aFFK6H1DXBbeLEOBknoY6VRnUNATBqTZEZaNaDezGn92i6J0ochAAjgZwL7VJ
YW9WD3OHCjcuDj3cog/qRDTtyq7jnlEkP9Lrf1hHSirPazF6V0la03luffgZ1IQMkzr3qbippVxU
H0c3nLA5cWLhVjI7vawNbJSf7iYhXF1EibzfNBgEoRwS8LBISODhjurb1iTrY066ZUMtl2kiNJQP
WzLCkISZBMQD3vYd1RAEwbIPxZlmnDffhVMlrJxV/4rNfKQNDkpNMcIKxF9+5ClJI21Gq+tgMcUw
ijfQAJIiwapkZeHXvs+67K+FAN8Tm58eSZie6oE0gij7KE5XW9lhuTUoRQWE7XjigWtdpD194YTD
bMgIG4Z63rJTydqpCa2YDH2XokwWdIeWvdpAuOuERQ/fR+O6tdBqKndDFxADobPHSXrOmrOLPejb
WiVb55cUwknhD9aJLE4EKSoWLabIVfSsSYzgrbdyjcUR5cWD2AuhEo5Q3FN+RXpkdd5Up/43gDZx
MQoHcdA6aV7xNjHm0fJo9Q8xbrBFgkFH9viZUPFcXea9h8GcTpJT/a5n9XN8IO0YYBTqGZvtPsdk
dGJipf0WAHiNnWCFGgz0CkjTasIDoJl6BD79zCV5BK0mJwb4ntObHCZK4R+/BSQzgCehRR8YekdO
KrX/rVyX4J5DY6nZyik9P1FtRgBbdhprEUY9fAjadizthXa9l6vsHZW7vE3MbGVhkqO7CRJkWnVo
0/9mkDdTr0HReQx1uTZI/18rPMcTVolraUnaQsMN4T4MAzJ7xBkLHS3fju9FjSyPVjI+GGSLfeqs
ZII/W+PY1IDtbKjDlsKjDlqhLlSSfmwsKBNq4CfyfGtBD6siUJ6ZXjKGO/8LDWoRJq1lJhVgRhuW
FhIdSdyb2oktl8nOottAbIWXZ4tEcT0JpQvP/jlfOp3FZ7fxQdro8px1+Ok8Z3IYIbYvQYPvP15E
sAG+0Ki8ZOhoRt1eG1NSkhqgwntW2pSyGP3t7XbBRfkScfh88S6VfW+O8omx8ZxYRHNDRNd2tPov
6DXJeIWKvJ6TLsIEcqZrs1jb+dkLysu3Ed+dUFSMZNlDgQsy0pJEMHKyXmqQZkUusV4qU5Rcmz0D
bBAdS9QdFSBGHqxM6XX9Yf6Whpjy3lv3pBDGImKyC3OUE3lKHEk8E95x2MBqwzBuUD5q72+jveZD
AFEEzZLG/ofXOY5If5ZYlu+HWSd8wnBZcP+DtUeCC0JXpsTdBgHEcXyJDYSPjUT2UTkg9J/+rVX3
XK620b0rix3vu90Ox2Gj2zNLf1Yl0BsrFTZJUWdMCu13STsYVCrjrfBRR8+g4XIGKkFmBrAgk7Jy
5Qwkf6qoQEsMyArp5O5PKzicwHza68xYF6EZqhVj+LGU4f361O13gWXdPGDmwvEtY6gnU1a54Sgc
43E+eDRF8ku2idUtUOBRs29RX1RNx8H9NTT/TvH6RfzbzwZhPl5GhsaIlQNbHi7KH15e2eKvjydm
FmJOS19WJqJFbkdRGjxH19Ttgod0YCwlgLHeB0qpuT2IeDsXFtyL0dfBYzKOOmQcBzB9Kg5w6mCI
9UUVzQge+aLAjsBdZV9zrHv4nTJ5rXA6pRue//EmmOVuWZyI/MiFBKYcTAVl0DOylhO5QXWEcPmW
sQYQoqE0az3Lvo1HjsQ38NIzX8lPr+ocIlzTCuJOek7dVFCv8+SMljL3qKhBDvJXr8fNm4vGembM
yk+pnMz3j/I36OTi6wpNbpZyltjYBvybPfer3951cJx0ZSnsocV2hxcUbPZ0KEQHWwNk8L7721Eb
Guhd2hjm6D1pOtK1mfSsylvkCPBn054MtaN53lZDYGXe200QxzCg07ipynLhwy1h2smIfY2ukXZj
bOG4+ULaG+P+qspYffUJW4VIYpxq7IGjSX5RkLRDcL9V2ZUQwNZ8AUASOzSLl/dGwKskS7eRUxRc
ubhBqwvh1QO81PrSlcYq/j7+BxJFxYZqFYW7uWveYw2tWV0QUL0tjTF/lPm/Dn5wdYCmNMrEjX1Q
QcbhLlRfpAsq1RJqp5K15a50AFOLrL9uoMzA+xsENVRtp69rG4IcR9/Dj2MDD/EuC4zTLzgbxJ1g
p92/Neq5+2pDX49usJ4lVvQQMx5iwVMmpyLZqVYPbZswdLqhiX6nXL95huTNoYIjL26dhlQR2ZVY
v5oW378DCdqsJ+9vt3jtCzQQWyhhq6QAjreFPFyhlV/xWaX284bY4yEEzjJ06K1LQ/XPPdZu1tg7
CPt61kezrEKQVxqHyqX0KCs/BPjdnzeWKb0i1cW8pvx2mEoANfjE+/WsjBB8sc/TpCDZgNz3CTGV
C3d5yDs9RBCUSmX3i2ZAZqI59/hC5lx0fNrewxuHBkUnKkyZlP+YwpbJh72bgEDTvtVHhPRFb4a1
sZR0IE2HaguRHj8K6O1spJTOk/vBas0U5VvdeNuQMEfhImDJNhSKyRVqBv+lS9BieQ0Ub5I8mISz
Z2faJyhmfU0FjKqyOF8OMcMcMRVTZuU3HkMZ/c27icJDPHBgu7D5b1qA4n/AwxRzjt5oXnMmKmyc
80utmfz8FsRmtdZapPi4frZJkXN+tuyW5+PT/5LPok1IP0+8OGhQauYmzZf/PnAqS6V9vSLAi43m
58uAllD9fBy77wt1XT00vcKoRqTfgLwdAYhho5tpkTWNEW2GY0r7wMpjMkRtVl52BgPjLbCFiPN7
g05TQTGB6NsNQYF9LGtrmjv440V982o/VFAHuMlRqZELIrsvcCNcy5Ee8ujps4afOn3D26jW678Y
FeID2a9o4vQRu46l24qteEfChRApNQ5Ctj7W3mzzQsKvJZ4zaHElJDHOz279C23Vtt69uvVUjLcD
jEDvLhg+cHhc1gJR1qtJMO5ctgl9zN72L041OezDcFiPv+xOZUofKLAyIhJP3mWUMEMAVRgQ5AiQ
PKg6yifh14jpPo2Buzw1eq0Mea2HY+C6NyhgFIVooBJ6+1gyIWOudCVWYhLKLWH1ZzEe5UyvbYBw
FMqc7k14kTmIBlrEwxq8GwK55L+uq9vWcAkPZ9Wz7pUCATWD9HlGTtIS/AOQi1U3URzCR57S6IFZ
H583+cROKmKmrr3wwCpyAtgweMUe5ghNXYhKHK03mGzx0LCGZB4F5G14AHie1kXGI61iJG3RD+mT
LoluW4G3VlN6v3gvp5BQf3AYACQWBPesRqtiRbIiNJ57bbx+oPsY8opql93txiAut5SBurm5Nx6p
T+0X5uIcVwCUFclJda2IIqsWD7iYW663OOjFuk0Em51qfNYDeJLrPW8MhSecQSYICTNJM2m+aVe1
EhxHMXx/QkzYcz7eIzazsN3/hfRhgV5QYF9pwhSD5aV+h1Nt8y7q9vPBS+7/zEHRDN9HUoCt9hX4
+fNHADzq4eszKk8eAEPOyc+7TTiRMM1fFJViwq/qtZJP1N2tYCwo5vhu1tCm7HLtscwp1K5+UYXL
ZkoK/IJf4I5dhLOtYg3MKZbTr3YHhbYR8d4+sILI6YkqFs5n/rSYLHp07B08l4DXeyYEVdotoCF2
P+ytjSoa1mMJo34GpngR/NetmvLR+bteGaTZXOpCHiZNP9K1Lx/ZVwuZxqUCb0RAHJ+rpVTyBVcu
M/eRes6IVDcvC9lYTVGD8UJ/f2/nenP0E1SJaeZIKplBZQMQVO+i2wwxTR6N/zHy7+MjM11aABIx
ZAhyZ2yrg1C51c6BMmik7GFQMaorHOpc83J7hIxXWflpq3gKqQMIVUtUtU7Cp6EaqoWmKHby8WsK
B5JLG2a7bmlUGRXNgJns11tE0C930pYlfCJmzQUqe366jzDK4Cr3eIvCuSDclmE4FWn1YNoxakMG
KvUaGwTjYDVCCQBK7ZPRAQBMLQgqod+3hwazQugL9s7zlwjmNH7o7JSzKtnc9VhDhkCiUINxlOsN
LTX56IYjxbT+2+XibvWBEpHfDxRsQ+XOnJ2pBfaSfhOL3Oc7uMODKQxOTCuPADKGSWK++smvE6bH
LvKWxQZG62mpMzhjPJhRmDbSnj6k7FJETePdOUa85IKgUepyBgS1UNsG9uicdbsZMGWs9+xdBCJQ
2fq2i2nn8c933iWFeFZW9NhYjgW1JJ5crXVZYQ5jRXL0wr9t8f15qxVupBWJQCnvbO6ICv3qJEuO
+z7LS7CteYO+TCdgNVeQtMxvZc5fiKzo0G3klbWx3ABbDuN22meQe1M0re83BXieZqirV4acPgCT
Z07LJ1CqTdflPndx81klmGrB/Q97uhoYXvykMe41J3ZvK3U8yOefhEQw3Bn6KMhFPZp9Kq+QVXRK
TxE07owLQZdbnOtJIodjAA1gDOby59VZUtHZN1oOKm2hCfcXoVCgn754imeCg70YI+iZShUAjyzP
jx6fW5Lca3PMdNxvbkJCqLI/IcoSnn5RBnPB+tAZzw5qLAVeylTCa9xdyaHcUsk4LaSD8jcFJh74
OyUjG9nq6WXee+1vZvNV6xsMFC5ebYwr8Ji4IMUOTpCVty/66kx4CWBKBAFzYCIfPSLqtSWgOtKZ
cM+Y/ax3rhpwLBmgx4AiQyPiElwuv7+YXTeGgrhvY2zI37o0BdKTzBuOY776UdU2BA381emO/cfZ
GEoBAJDhVzXKnmD7S7PMlXk06ATa3DHqL5/4gfd0VBB0bQgt2ZtokG4PKDfezH4HW9H91pULjy1s
zDvJ1oIZqHU9ONiyZuISZi93q/zry5nPqiewV+w+UNOuWTJtS/8oRTgbOmGKzSJ3KTYL335J9IFo
DePv+zPmWVWmhPKAiFIQnT+ak7Q/I2Q26OLUGtje3PkEglbFrGWNPRqOl/6QbsfUowmPe2Zmxpth
EJrUwT2FOFmIGKuGisPaLGYZQDy247Ck/H+2XiXxcechqwDqjd0fImH57K1xvRykwFccyzktkHCx
5MZqTHxefQKqaalFiT1AqzQGUrRarrzdZtFxGLRzYn7Wpg3ycsUa7DunSf00cXUjX3lbL4vV6nc/
LGZIYNCy2bAiXWnjhuu5nD3FGCdsHGUK3lLKzq+CR4WY5KW1PnqNnzsBa4vlKoCDBv8w5yojzZrK
Xlx4FTAdEg1dAT2iMolWcXvlE7gYMqtk8uII6dKIa0Re/InYEQwWMELf7Say3NfzEP4El4dskreG
23wBDVki5akc2hzYytfd9gf0XvgT07OuuGoK0IYbmSqYdpbsYc4TOAdLGjOGBeNvH/k6c7n5b5w+
f0y9h+4l8y/lGH2x3hwWXqcUzphKLMlZIBb5fep0KMsJfesgPUTf5ZJnj7NQD6ReD/se78wIarLz
thOBYLR3CnpIvCKbBfonxXPVr0BO9zOW6buKH/NythYFCTJRLINTgRvDiUR1uzmUq0jF3Cey+sXN
xzmHanbkEF6s6u9ZsBvcggmcb0YBpCXBX1FR3iyavDMejHmPUROpCWBOZmG7Tgks6PjFyaG16Uz5
sEyjqjuHdM7vw+XGQtdzcZlW8TyZpQ17BVp/ffbpNdet4W49GVuwd302sPUD8AiU++1zYTlsfP1d
aePaaIKUcaHqotXRXinZHPHBTpVlveQWon6fNSbYvwiQkTxA0Fi5wNktMWQz2bOnehh8g+DGwpcu
drHey7L9odcB1xVOLAHYAm44gy0BkFXqacP+m+wEuhflMc23igdk2MCQ2nhU28NNfcktw6QyuqE5
XqdFAZECPnx4b1nB4pkO5ON+i5UDdn1UBRGTT7YBQKza9hFdYZX2b/5YRmTJKLtsKBPG9MgeUCtY
Q2KyufONdorO0Mo7UtokltCOxaWcQB34Cx9O07FsacLUMG8PCnyd3xTeW3bapuR5Jgnep90iAmta
Oe4Nbxc+5SbWBO+j6P1n9jmE+VHK2PzKF3oUwwU+ptY0CgALZqRqRZSmajW6E6IjeVo2gGAte7UK
TTY3FThIvbI6OtoGaOtQNAF/7jaVgc63O7xkbRbv0l+ZE02dkY6q3wf3pYRLj/GZkJGPI39auTc0
apKy9ohZA0mtBmMDJ3e1BtNhZoP9ZRDfw5ngPH7OYQjF2I/zmQqzswLPgKCvhPWmBOGkaDVeAcI5
T6SMto/+/ApnPrlfhi07SVWpJGnCNiCt404rippkBkzd3ag+yjtmJljd/NT7zNngKRUNtY6H+Orj
XrvWJFD7AVQjPm2gCulWlBo3UiROi0UmLVBLgdPT0YmObVofawPxQDWZ8GyBHSqvyk3CpLAj/Ajj
zUfzYseayZt+6LE3aVXfBt6xwDX+uFc1v6KxpD87R0MgO4TjgkWo27dJTp6v4izI5zc6dtuEQw3h
pmKf/fnEYx47Ut7PjcH9ygqEgCXeEOVUt+/RyAdR2BMytmQNo4CGpTpgN9Ts//5nQaC5P+a5Hmby
7yaXSqvWdehsrZzPjX1XF8sYPbo4Kr5QL2zHT9KHG68mRpXHHPKrgC3PxY1PxdBFvoaSDuSNJPEo
ZZNeVmO6sOo2PQcom7TbgD8DW4Wz86DbXSRV485dztFfqSqRPfQ0+Vk/xRjVaD5wdbTZdlt3t7Fy
XJjw5zjVcLY+OscsmQYKmPVm/Xpwm2ZXIgkiiyJiUmToWHHMXPKNfQrKg3viHNDhCOxVqog/oxoS
MUz/WVI0xQXi1WiCWgTXy/vnZMf2qb3CW6wm31ry8q0uc/4/l7NE4kAQupt77YMZvt3VPurqp/BQ
+fg5zGXfEYT0EurDhAaP6lqzuxjHIwlMXdT0TyOSFG6/bJAdh3VfXgShCpkCsx36scDJxDzEOYYb
Qc8jCWzLg5VVDnLHaBxl95EtOc+cwtz5vWLhvQRlLL6Ta5AygCjX8cNWUT51j4+cP/jk3zYfjbSF
HkDRYzWRBNMpVL60OU/AusvbDOQ37oGToGKLdn/RHKwESiwRpcozSIhKBw5YbxdbdN7oKurLMCCT
0nPo0/YAet4bPKvlAHG0U4D/uzwDdb4kgZWbgJAyfccHXic80uU7Z3MTnwpgsgyG19jjM+KXbAR1
FuJodWZcKdivXTsFDisSHYF6TC/dgSRl/ax2HPMICXdt03WEzun6trMHCqqkzPiE+L/mPHCisNsL
QnqDh7i7Jkk87oyDPoWMy4IHQ/qPOjAZJP1/VNC/5pMVLfcYLX1SPr9cZoWaVnxksbYnQxph938p
k28Y1e7vHwh/JCT06sb6NcPZHxTi1bA/nq7dqa9JdDNNUCTM9jwWfq4EW1Dv9uUT9vHMb9HXc9IF
QD4eIQZypk6Cp/UEdGuyYBBbB54/lDmEAfLRXCrZBNtRuOMnStSsitzWgyB6zwaIBzbCBKneUx4b
betF61h92FfgjL61hS7A584o0Tlwqp55Xu+7+94ONeJn0dOZaBVG9wK8M7viNh3m1Eng/1Yyxl0A
r3Y+RswIL9qPpAP6pP69aBtaePIzQF45WOujBa53I40tP+J2dvOxfuwrePNB9+DsbeIWaxXChQRq
9G1N5Nrh1n5rDU5h5qweCMW4ZfsyXa4xDTbzzCW1Ee3gCZw9nwXT+Q0fqqEv5yNNgEkoWRtdkV/7
/uev1PCLlzscjLW4nwXVWDZpe2WSdrsF0nvjN6EXnDXh/bH7uXz/MqJ1NomnMMePGMCwsVMP11Ax
rDPJXWDXr5uB1BNxDuZi0ADrZSgF372r3fCWvcH4gTnsFXn6Mn1SPL2/AZc3gKs+5ALSMOGX2QYk
oS7Mt241rFTgvV4Zj+I+IWf2YziBaUoybGMVTfLHpY7s1jMcL89aTvY8IM3x8rmNOcm5OVDyvawr
7uBPKYLdCKMtW6zIbwMiJVIj4tH4QsnnaO6Brb8B6Fxl3rq4CuNwACs/q+toBOWB5T6dpyTyRcLP
HqHAvt+IxremfJwuKCzaazqKQLZvfA33IevJQjdVNXdGw5Pzgx+0c7D8EGdR36ourZKj/jvH6Vc+
DL4uVwgkpRpYEh/NZqLl0ineWqbf9z5Xv6orcEeT5ejQC03b2h8P8YvXTeOSqZqf3ITW0zpZdPnw
FWyUQ/WhqFnHJsspgK2BPJA1vRfXQk/E9FyT9Sr2hUGhIuRAbLcX3x4mkOoz/DmwsqKWUdLQnsXl
DwP0hzl6Uzk8+2eeG5VTTc0zuLzUFCYKc9VRlqguF5w+4oZZaPmlEbmC6yQLpF4DS5/AGOTFcnby
39Kw4+63gl/HgJX0yYBuTrxh5zSulVRGrwCwLwORvWVvnOLbhLUdNpNkuirDJ+LnrsmHBnqgLpUM
QEnpofDBvZc2gf4H0tnsc7FqKW7cFAiqInR9heMFBjUeeJ5M8boa7s6CWOleIWAd4Zd976CCp8bs
zpDosF9AwX79XJ6WDaHRT+JVqQSRUKE4DkrQQoImhudQKG6hJS8V9vB3dxGAPaVgGBxs1pNxPpiA
GF3aecp6v/unCv8TX6UIDaccsj6gwJKBSfjnsuDNzrXAAPGU2bZtAbYScLWE1RvWcL6Pqm+K7UPo
8bi0AJ+uUlK34yADmMYJIhySXNuNHbAQBDa1dwAirqxnFwYTkfMWyOgiCP+xQpmopB9d+FNRI4O0
2Lb8JGfzsfvSlBO5NHSMfyhdQV7VZIcbfmoeXllxBk7nacam4jGGLYYv7C8jPldNb8HlnUvopVOT
4gGYj5Ic7lZHIKjHg7qga7vE43KoTNRgAvL69R1pt/vzGbz97w5L6HYZv0tCwjzoYSiPPkx10Xor
AQ5jcIyzMUgC3eXFVN9pBvO7zZ6INfZFAPCsPcdsfbeO0L//DmTxgipQzo1EPUWuHYDUYppGUpmq
3/HBdLnHfq1Q+VOG4S5X2/Jp0IDa0hjFN+Jrh3+DJ437adRor8GjPtiSbJ3JRP0hl/sB29tDOP/s
JtqhqTv/jw48AyghJ17gvbis/fnp4Ox+Z44MsWbpbvAwluh/wi0Nut0b9jG9vVWKKLLKq9Nh6ADs
B3TOLreQdesFlYm0o0mTovegoWxw4KmqxybMff8c5gela0vpFgQCydB9YfnbFwwNV/vwpdCvdHGF
4wdqe7rUttNfW0j+tr8kyZy/l+tZeOMuCpEY+4HRyBSuAw3p29cQGVFv7/8M1fDKk/uFcBF0mdEI
FFFeVV3GDRh5ZuQW/FFFiNyUFih93A66VX8ZHCTk7662yKCzULcyWawFGfA4UEqX07ZnmMERm92H
r7koW5TNIXXW7PhRPZvKxYVleOBxyTfygwYFZsqRU+4UM/YoMMOJKA5VDqiy4n3Eal1YJm8/dZa9
G7yNu0x5Gaz8sA4MH1mZJEQdnVJmsgYLZzWtIGYaJMv7O/NAvBhFQueqmbQ54WYfjeR4xyHvpcJh
qDV0z9wMNhX77RSaTQ73YdJtQZK9KI978mub/yCU1OltuCwCcCpBGmodnruoajmQW/iCmnMWFNNr
wdaDHXF+W9iwZFBKWUPvlS3Sc6+bBkBwD2wokoXb353fN5f/724TSw+N/6xhuvhM9NfVWFTFpqkz
BloEuqPLL8X3eTWwasMEsQehL5GyvLUWH85s/O7Cc29CwZBSdGW2J5wasd+u4AHhFlgwN4ApRZuS
kJNd6baqQMcTjP7NHDnm4HbxVtoOpJZ2wc0ItMSngk/eknmLjJ1EfOOkz2nG80pEUrlIPUU7VrdM
WsGptJA9bIXRs2HI9JlwkOtvzUFd2ndFmwVB9OS6J9Nc097ho9UBvcp4S1dtfbikio1ixm3sKPw0
tDzmPHvOzRYmZWK1VBt5do3NCUmp0yWx4/hCLdtP832CIE4rTv18f1knTz+RvUIvsHquttpi77FP
Ud/10NXkhNW2DGGtKDqEgyGYALDXkvr0hj5DQXcfrRpsqsEnhawWm1GedTLlVnoTG4lAvTy3lQQT
9MH+zOOKmDTcLcAWRR9iBhB5KH14bFmfGxSxdUuHl2UDrZvsKUQzoQtAH/zyt4fyhJ2shxQItZIN
PW3E4EHmWk6O+0Gc/+C1ViiCwFdCTaMcoE/ws7NNBDfFo/1fceEUIooD8YcbRbBPcfEhjwOVxIdC
QNQA9WAUZlbzlZEKKOhyPWKLrCNaXKM1t3iTbxQux4ARqTmOFddRbGwDo2sp9pE7kME1Ot1xk84I
P7NE582/65SFc30EJx0VNn2ilW+ENC8W1OvKWxAnihbDxSU8Kz94mHLvtNb6DmlCyU3B5jcJf/Qi
16iSPjhL0QgL3Be0PXLja+LGHmPOgyrSBn6UtMe8GvWVzF3KCkj8BJ1+VFUEM1KP4jQFGWkqhbpW
7/XwUJVOkxGAFiPSfzFxahddLFkBNNsrWKwJp8rw9SkBreFTukpGb6kaZ5K4C3K+QsVN2fGzkcfj
+YwEfl7tnLwD0zui2GeOW8UGRToC9LXzp7J00vK5MZEP99W2pBuyKfBK5D5JS25h20mucIu6IXiX
IZRO6CdsbCPHSpkDdloQVq84zjEHzD97YmS352TkGpitIc/ULNYF0Q/TjQqiqimldUaEWO5364hF
i1XoehHY7trwIKPVyRXbD7//s4ySpGGH614P6f4NEMu/uVOQzCVqWYljPixtZEaxMpkvbnFbR1ZM
NNMwPGzt8kB34ARl9rbPPA/MDK0gP3wqHL1qIpNMtj3qhMnoNvDEsxdzpiLOIoVRwdNrDM9snfF8
8kuSHaO3Yt+0lhMDNerpwa50wL+AeABkfKjVBQMrrYLUxn+5O3/rkKSJLpOuaiLte71yEt8ElhyU
gD/fSIK9Bi8DFHYDjuFpJuYSqBwKyA6+PHuDWr9GNVcjx1o0wPfGQOGGqG8q8dgoU12LWGXJCC3r
CIkX6aUMG3/66S+YqpJi2CPDD7IrhW5d2cVufhQLx9HUIFh018R76xMLd9ww8laF0WgbIeit1pVG
cFEUk4m1oOHkUbP2GWC7gHcyTLlROdjx+MhLktkVWzbwhhsMre5pqgtyg3qciWhtU6wQcXGJlDIT
AQtJcZ/rbG5dsBPWZKJ29duBXjjhLPgJDAZuG5aZ+sY9o21n5SWg8ewY4xQIlaVOI8lwoV0o+ahQ
2ouFwQqj6OtfJhoo0hz6N5J9SdhdAkcgZYwef+g5O1MNzcf0Z81qqGKO64HubYwvPC11dgdgcn6S
3VR6U7a3rvU4pGFLrcy6YHnNYuoNMXIxakYucuK0smUDiH1zQnHsa7OKtNA+SUSZTR3CIpoumfaI
jEj8V58nN4mrVcciysm2XZbX3pHY8iERJprmnPn6bD3U4LRqJYcSXofTWgb2FTMgLRFJdbVFlot1
IsTnTUwgp5XBnk/qUWl84TLRHBcq8VjOPJemA1R5ebUEZO0dar4xfPMXQYCakuK22aFkYg9p6mpp
efSVB4xUeg+EuGB88oCD5Py/6WVeM/EHMC6l8K+o+34N2u4bkuYIIUcsajGd6YBkmJUbYRdpIHTN
ggW3X3Yi38sWrg1ErjoGJZmY+3X8pYOLoJoyqPauaHu7XCBPByTpPr3nkzXYJPhWGLcKmsg+AKZK
XUJWTK71jBHckGbv2HJQ+UqW+G3AKgTm9CwnXjhQoRhujZchW6RgmLejBJL2FcfttQ8Ffa1IUpri
XgAKb8xB0zCKjgRtomq41YU8yq7N/VW5PAb2X+phLx3zGTXT/ZAtLvk3mIMj33QZa7aLc4DIUJ9m
9nKTHZc3v+W/JtIWSynz/oUB+EFfudSmZxJDOrcAt7q7vHYFYdO4hoIABYBqeLfHq8GGzKAqeG56
1OboZ2GHpiMVIokJwcG5F1fv/iYjKumyODhMzesAoAQACWgXd88Lc//RVpK1JG+LBfdWKukRJnfq
1NA7k3+zR2wVQbUHEUHY751VErozfwShT4V7YjS94Df4RnXNBKn0wrFb35+csf9ndt7ZPVIh92fB
d02eGR1o51YP9lORlabZ+jBB+ODD/0uOxkGnmR0CVAtywtyIJh9ND6Z4q60HaAUtJVBcbILzE9qA
5Bv2zlKFjJDmfW2hMNKK4FIdS5cQVZk7IAXzAA7oy2OBS9xwgTwbu0n3bUjpAwSRbgJuDykF9QyJ
6tOhZ4ed+4NWNRT79Vp1dEE42boiJjgYbV1FiSIzmhE3U0m1dgPLYGfKKxJWmNIfvKePn0ITIwMB
DF+DJx/QUnIXaKfG51hnMRtuuHkD4XRQ2n65PvfRtZoVmH9b/0v2f44P9HZk4jzb6XH5gyQAy1pd
bS/yv//SfSJ3ZTUOwBUiGYafhdGv3GCcBlJWQZEi2inAEGym0Ob2BCcbETp8SRlMJJx3sEVve4uu
K1+VtTX5RNo0Gn1sSDZKoi6yC54qmzkw2N9JZhcWrcskP/EMUm0rPiwJ96lTjvJD28vUm5kC0CVq
n4vLVPUyqG6n4RHvhLkgSBizKyT4PfE9WYtHcIE+KL5VAnNYA6kSOMIeXo9x9ejt0pk/WcTyTIHa
ZHWb1p3Tvyj1eb6C+ABDomHo7DqT/z7+dMLSpJdDrax4ynqP+MaIXZGu1A/yMxNhFFuOXApZyiOy
1YBk7Vf5PhQJNW81Y2pqcmYyLoEMDt5prLs99MH+093NhhH/FNbxVnzX9p1vY0JT4CRTxJ1ay686
JH7QeOmtS+j4uc4yVPLTEAlgUkEgCrkz0ekgX+Fcp7ppMIObp0G2Zh/ARAQagqQpWu3ThqDdmnPk
U0Hsv3Ey2hbI5b0JVGhTiyAUBJiLwlS82MxXkxA2U4w2g38kdtAtr359f0Cbw1FycsAAbseHXIr0
I6yE2+o/1xAWzTe3d6Q+nzGdQXyK20i02qPQZHEm6pSiAcAXxnA3LtlOzgb70+K5N+RqbpbPFpKV
XA5TihRTqfDzYr2bU6cfELFn2ePZlsa+nfAUosk0zMLolKigSoP2cjd/89AxCKZg6h2RHRUnmGAP
trrsshIxA0OUFdWLRhMO9KxdnIetF5wRV+/AMmv7d0cArVBrQmf9dXEdzQAWvua/RbX1fjCvyuD7
5BICuIWFu0TSB4+kVBo2f1XDuP1TWcuSz2mmE0nXYzqLx60TowRlPKZHy3TDzYG/S5RbwJRlq8iV
ra0Uan/rHD3t3UmUCr/GBn4DCP0mS50blIyEjB4kubNAHqzm8nLhRJ3PUrLwF9z4gv3dXJLNG61x
pW13UfBMurXqOOJuOuoRXH51JrNBzpRj5LoQbWykFZrTwRvyoLyysE8DkyUYYYyddkugN8DrLeUc
qXoirCbHrnFaCdohOwYNt/UBMdxomidaK4te1C201U/mckW8B6h6iNxqPeNCJT5reNfrATgNcAKd
4eKiQOWKQDOBb0KDeOsfyghkGDK/qieOw8ZgVY2LPfFqfIoVF0WTTNUX5/LOsGTfe4RqsteeL4Fx
70ynu5LRdrkl/0xkujSAxaWIJ1NalMUJCGK9wuxJbqqqhUauktCGcwSQ+ykyul3iaRVb0LEB8Tra
REArbcYykHqkidsyI2or4EqVcvgfSvyhoY2c13TGvoewTvgexrbp9vlH7jo9PTvlt261jWYoG+fJ
rOoziyKxWw6c65sgnCP5ttclViuy6MfzMduyQukoJ2VamloCgEwmKZA8MqdUZwbNJMXbBkzXaXew
ZeOtmQfgqaoSCosyqPOU+n+17FJ3QKTpOnFJN5UsepmT/YAqicakRv8ZyKY/RDx25M+VzVDm2A9b
2NxtpvJYOqA3tVQp67/Nw/uM/u1DGKaUQl7lWMjjcFwT0IHmMCFJydUPxBMlJW8/gpYbr+GSpTEw
ihxiVu7fAR8CKjt2kgDrKi9Qt8ZkPI8C6gl7OvuQxbg/zs/nGSTU4XC/sBTgu7s0am+qnas0hhjG
x43ii15+oOScuXHDLP8fu8wA+Vm5qQcQ7W58jecCXYIHDqbvLozAIhpHjmvogu0TRSMALNBRk6bX
xQRlAnYb86Sqaj/zVsKqP/xjB5ChwiXt1djW4fQLoX6hmKbePxBefLcd6BYJ8heUoQ7UJ8BlB63U
OgsdcMfxdBN6B6zp57o0HVJOqZ9bBK7H5TtBzlXiBoUQ/fARKslfg/5h6yX3abe8wLH60HRHr2CA
KSJ7RGjmr+ZG62sn73LJMh8tPOO9a4VitBC5I86Kzu4yDirJxCZ7oTfdf5ec5SXqqUkHE4fkImLz
+KJjoZjK0zeTozD0CiRxmiSgJ4u9xAtJqhSeWCNjWEjgzGluRCQVPlCJinNskISU8LwQJALbRsDd
8YJzk7zcZPpG6hxdeUNIMDCg/nkt3YUTsoEprX37LmFnhPFcNuP0739XF+jTh42EAExi/vHaKrjR
hqcTPgXV4QrMXAKPI5BqNgcWzznk/oip9yqWMUHHoSWCGTLkOHPZ9ja4XKkyZhCrhnOE2fZ+ERuO
IXv1HzqHywsXVREcVgRAEM4YLgyqbYhgsu0UVyhb8ShtKFesPBU+UVUjSGZMbazOyZBBhRFcp+LM
bicAfKf4nclNP+HNPeMVxP49YGlx8s/LNxzzu8pFQd6L5tyPmQc07jFuauFWUmoFzeX44+xb3uHk
giXci7Fh4ZiRLxwgsyKZfJyq0FSe2XO8eGWa5VKnYvF4MsT1cCoU0tcujb7NjSLyCJccSzAkKTnR
ojgd4AboauEfryot52Kha9ebZLPsHZ0zMz6oOqFhV0PFSOQb8feba3OoWmAezoWbT6gSe7FuZ3Sc
bNVDr4i8Fnb8BJjKclqH8zU0LIqLkmg8dA2WN0je7Sv1E6D9Z9j3t4IAc1DjQA7afT7TUzIxaSW8
evxEclTKBoshdW9IDIskJATYwve8WyYgRRbsKtPQ7JiRI9TKe61/l3ke5CLRNXR9J2fwHT/cd1Df
kzNQ273d+QwjOo9P/vCj3UmZoO8JEjma5z8PusXmON2jG5VG/RMr1QvWH/jFiKLQS9qR8E4fjtQm
QvLgWaOvSG1HvpgSIZUULtC5E20olrFtMYYK5i/QczzINqzjfwb+vfNyZovJEHwB39du+DUiE32I
yR1X/6wwToWn6lxCTIGDyxDFhfvUc3hSe2aGvNz5LcVxLo//3XKnaCQ6ogkH0jzc/sKYUvJYPyLx
1dW5hI0iNFkUDyLP85Pl8W/28qGzaF2HxGVRCDwn6COa8DDtD/gtmroHjpVV8tyYzS/CAzXRA1/D
lpGk+ZUWUdIhd5qtiCV6QthiCNtKhuRs6fT2h5idlOkqzqVmOiFSMQ179AFKIoFfvaDn5uLEajZ1
47mxOWVeJypbOIwFP/dX7Szz7KqYPP6e+Fo1hkUlVahNgvhzfiq+j9707WnQu1aHjX7qmTLq9j3L
z6Hc8wcytSAmhmd/Gl2bgr63lQ0EX+A7nD6DvfgLaGZLf/mY4Uu4rDIKrgFXA4+lGz1MLx/Ji+Z9
Ui67BxBP0bkiYqD3qF3tgOj+XHgfMRmSPYZXPJ1tw4RUowZiGycHesA+zl1dYUuHTbwoDAKXaHd7
K9ogsqfbAStPWIYULZy45Jtfq2ySy+6WAGOnINLW18xPqszyXi2fXRoHm59awvhIC+peVwcmpJwC
twHr4whrMSwHlgQolOeyCd4QhuWrJMpndHcEENnYIif27FFVLRNgiGfef7L+hoI2ER/uZku6LrmB
lYKMgG9kINLvKwtCUxASnqWyzDULpjjAaS/F4bPJo/Zn2Z/HbBnW6QFV/7E43ljc1IwuXyf5s6Xw
zY/jdGKD3+KXlo+H0Mn7ls38u3xm6j6NrSETZ2bZ8Tl4shsxHXJRsZtzuaKi9ohZ49L3VJ+xje8y
BYUJj489shJxsLEt2OqPHyvO5nFNWwedtqfzrb84L1jB1HwskSnBgT5ecI0FuJEH0bRgqgpy6fqZ
UVLb5dfCUTUDMmt/EDSxowOTCx6iOalSqfAsC6u8lD9gNvoUhkRrnCo1XBjmMKyQwQjybRMvVgCO
M14RRxZGYO+JnWTz2y4IqJP88LYbJNdRCAM4iGk+bJUZAmj7Bvocqco5siqNPF8SVz+VHaWQ5Gmw
DRqjfIw5EklDhiM14t+B0bqb23FeApHdWz0ELPmJp0C+yvKpWQwwVzDVOcIsywdqEUYAbxqbqXDh
XHjHvwhFa0gXisNHFldcXe6HZpECyPUZBEKHoXgjwigNQoGcC7j0Z82L9tDzf/Wt11DA8tiXfDIf
2KO0eMajd/8TODNw8lwIE/lfvnPHN5GFg1WB59GbN68KBE0x56N2OCDgCpSGp8duQImmkS/D4tFp
b3NQrkGIAoqQN6+tPMAQqfDIzuDkm+Hv+mIEyEDgUWFYmnI0LO6oMzYo2C1NxR1Qg0QttLf6kdA8
UbSPrnrNXTLsUwSKsOSMrPXBegk9EWrFfY7fw/bNhc/xzz2hMyqHPT4h0t7u7/gmXRe+Io4q+HH+
IN23HMm7T/8Voiul/tZZ0O5iUboDX18KRKkTU0b8m8vTKJgL9fPuril8egAl7jJbTZVy5l8twHAD
XfWWeob8u6Y4++JsB45q2j+t26uFOoyxxA4gXDpT6uXNwYfrR7QZ2z9Ug7ZiLSAcmOCP9ibQLmoQ
0X54983SnxW9sCUNvv8U1WYq5+lKl+70H89hDCHx0BFUx0sRRBQGMLmTVNRclgISNBjnP448+864
pHteDEqpSUpDgXNFBdDsjy6dvD782+bl2VqSrMKv5ByF1M8iyGHfD3iSk1VKYp5t9GZw58oOmF5H
bguq2c5d3oY5ewGwEtw/jdawWSUzwuWAC7ImnZCZk7ULXN6dnaXJGHwke212L9B3Pbs/eUOUk3hg
P0CWvkU7uelferV1MqRXQh8ZeCpyZVIxUWk/J4QiwH9+G3QmvY82XLLg4yv3Gpj7C1nrDfSFLGCB
plg0N7uIIp3e39L+AyNz6B284MuuZAYY69Q9p7yFyvmWxtAEf7odvpIit9HkEvk1xJ2XPljcCbnK
vOoDQ2nbburG5QL+mhCqAsd5Txv7ZscxZU4vQ+JIMPSP4hIgJ3qUj07gr3ZbLfLvpvQo1A/RBQ81
SVbb6MxJa+J44BkOrKHWZowqtKdJ4VWXTzhCa5FA4+QPwV+XUPKFb0cxsY8b7vuvqG3k2HqFIyu9
WxhyZQnGY+46RdXO9p0BZoucj+KRX9WRNvQrKa50hy1zoJBj6v+k1euvGZQHyhXBPYLWulNoTvKc
S1a8BwcY3ZIe+dxiM3te9P44xQQcju7dTGLKLR9xN/qBIrGSyyxgQCwD4MBqd2zEt8md3Gr0TJ2q
004Tzgb2SAIuAp6xHg7pjQW6flTbf7JgqVQynVz/GghMHd8iHwU0QRioeOXSQuXOqfhg64LWtI4H
Se3QDP6Zb+aLs/7g9ma46t1QiS7UM3edDmUIorPoRCOQFymAGITCk7fpnPhAVpTG5+FjsXf2I0pi
1bo0CLDQEFoJ9g+JZw6dWcM3FmvidF4YdI3bUV93It+azTv5VRBBK4oBt/NEdNxh20fi3Knbtfia
wWcYQP9bFPgy4bGR85A0Ql37qBRMPdzHJ2eZmpJf/MzrAM2uOznwCkUyfCTMFBzgpp0SyTqZLYzb
OKtemINQ8GEoSBU9jUCXmFi8NpVEUZ7EDRJfCAtfZqIIxMunUdpHDk5W/Hie67WtH4+z755vS4Zs
T4GebrRSHeENw/OG9DLrEEHYxpvtf6TL4VzBnOo4SWcQxbfs5gve2EGwwttJJMYC2YTIJRwSbZpJ
Wugvw/cNi5Y+R5DtGwQ2jAC2jcrDYx2oHN4Z54a2SC3YS5bVsZClFsNlYMfiGkECM+wbA4JuFYvZ
9tpfY0g6IOGm6noki+NfMmEGRsWm9ioDCZvH1q6pzGHms/NwFUMXN9cYU30A330yRm9nSnRAhSAW
OipaYYo2bt9IcYhLfXZuTObs5ohIAn/DueGqaHuY7JEfIFaLWen9uTRPbMohdaWTOseiL6J5t0d3
ztZ++xnR4SxhU1zbDgK1lNV+XjNMcCCkuOPPSbpRGf7CPQIOgLmCabUQgVrEhliUMey+a54HKRzL
ZxKRjerlhZaZcBlWHC4MgeLwR4pEnAyiXwbVp9grDvDDIx72PraSCRNQxGT3V9K7JO3Eejy2jyk+
kAsGmLNSb6xCxRkAcoP5+AaoSuRFhJZ/DG2XWK5+AxXkKPjlKruT9QVrS4l8xcMdZus/jH6ANyBd
TkbNLpEx6uLvGxY0htIExm0vb4MgyYF1RKZ6Ve54xKe9An1MLUfurbmgQRDUb/f46rEpV+Jlcp5L
2xhm9lyhw+JbqYKxASTAmDFz7BN6llD71CJ+56UyVKSFM/ueDjaS7Jb0DCET/eQh6rjkKEIkYQoS
NplBG1Jfz1Hdo+U+paV7ia36EfAr1ZHoo9wojIHKIB0HV7l2QDPGZKYEbwN0The+8AkBMti6Kxm1
xBKYStzePDO0pEPuB7SRMFw77zXSVtiLzlTZgJerccYdgnbNDPc2s6rt7cXko9SPaAhdc54jHszk
BxcdIdFgZ8c1LDj0wtPgZrgCD5twFs9UbNUY9OiAOyOJxx6JQTgRhAmrpIFuHH2LKjz9zHKDVqyP
mgbLKKup5SNReVfx8fEhiqWGrkrPsaCs/2tI7bDTOBECoOsUInYns2bwjdNn+ektYduO5I6etytA
4s1kB2eQH6idsjZfn+g62RnUrEiw9ik646GalZiKyce+YzF+/VZfi3bsvpyXj/Dumwxn5VZXDx0f
4INOIk5oYiWKrePHNOR9aB4+Q4cVVIzOuOTSnnVNNCgPk5rTI2xmFRiGm7rV6uCAYVYLH/W9r6uD
8YajEpMMOPtxsnSwSo2dILjjmVqamOEgjh0OSaWcy1+44sol/nGWy1/DHFSdGEt4KkiMa0Twe439
4m39l4yOIoNUjmgtG9RMLg+7Uv+IQyPVhs+/8rB50d/0n2K+Pjq6CCkQUi3Tbk7BONZrGtAm59+J
ngN/AQi77MfMl8DMb2poZZVia1tjDL09ntW5boxcfvRSp12PH5CRBofLG+yY0l9z2vKTHRyNhehh
/qru9L9Qo5SvA8ThOgUc4C8VfC1G4ZGZYoYmIVtGI5HXgScwSUpfPN1AQTXzYK7qwMV75q41LhC5
oCxGMEgbrBvvpiZTDSHfcMnhB0JLSQB2x3aIzZTspgimCBVLvqMgqJ23fWB6ec9a/4+jsT7Jui7f
8tieti6lboRk+QFti6Zo3mm/lr7ybVtmGq7lPY/MXt4KIZ2yTFtcOemXMJQeQvf9aAqLD6HmxCRN
xh7cOgfXKcDMb513g2zHIVv3B0bah8xoLqISPGJU7HdiIdn+M8AYbJLZLjqXBKJkoJEe5vI9wLRz
DdsTD/EmGBrK1vrtbGgNSwWN5Ev00DDYdecpH4bxum0I2tSDOaquAK+mARkFmTv73OQ4QpGqiFtL
UROpqW5KVRluHL6EOry1AM1tH1X6UyWVCkFpV/Cqsoedl03cmRM2b8Nd+3AQYTJAAMS79En7faIl
yAzZjAMcRz+tDC4JUCWnCgSRns8LwLK06jmVE0hIMhgu11Z5ON+xyXA4xUCLA34fO1j7b+NgnFoU
xQ6BSoT0/6aQdxyOTfYOqW2uD0aOC8e0UCqH4EvI33xYxcrkbEiG8Ch3zwOZmsjAjW/07F9aBeEC
cCYbMNrP90/oobKqgrHiaIfPceeldKrQbHupGsD/wYnt+go8/UrDA3lem/6V3D6PWmau0wYN9j9w
ruI1TIDRBvLFZBznXdcKnREbfbCL2A791E8RirOFNYJUNKSEThx1I5U/u2rA3xHg/bJMRmciyrE3
z8Py2UMC+oMBf9UduAJncDXg2IdaTXsEu4XE+zn84td7wBUdjksB5yADO9vB+LNyk5cZxgeolOlx
7mT0X6yFiWldMKMFMCGdXvc1gFQrYNYYaCvyDXW5126RgRGsscYe6qQ6OMxrsoyUb7AfTFK+VzKb
e7bi9eWuIlDNiobXitCePB3kztQr07CdRpX2pd08zw277YriwQ+yGkjp6URwnC/L5fnoWlQwnQgk
SBSXO21q0MMYmLHEMOeZrLHeOF8M0phBNqWoB5ezOaoL4++GMAVnhDvsZ27Boh0nFBEYQiRuF2RU
jd4778JjWP5VcWsMcz0MmU6bO+PaZX6J3/x4Lg6Lr54MKfPJt58J8VUfrSVT8TxIwztz2ZMo5pmz
oQX2VJcvSYBSjcF0z1J39R9yRx6ye/mJXwWyr1jbzizixOMiGO8y6T94HFYkndK9trykKdrzVpiX
4fnrTEnUKUdpEgFgo/35Ox/wvk7+cfYG2e7stbsaygNVWC3eMOlq8aE84Y0UD11ENZW+JAXLcipU
lj5Gx5b7uGBThycQFsOGgTblPhVaOJ6C+4xpqZ3Xcva+A5R1NkNw8e71AWpr/GF9mQf4IWCIQTLH
lzfBtN8a8ZEEtBiZmZU5RqtGIBs1ap/OWEne8LpTi+EYsMlKlr92cuMTvmrUXL6nrJgsJIqUw7eG
W2ow8mgutwcSLzIayI7uynjjuvmcd5WQyg6ECje2qZ1p2GKo9aWuaDN10FRe2sD9iVnpEjFKlOym
/Sr0Pto9IG8hZPJA220VcVod+JwItrVODUhOL40AplUxjcbeX5LiXotBkUqK4ar3PHRHq8OtL1HN
Zuk1gRPV6BxUmEjH8v/T48U35zoXByicvM13qPaSxAEn2+EHtj+kIqtAtFWDwFZCr2MHG3BwDxi7
nUsYD4xQubDtKU1n6y8F3/npsncXADlBLrD6F0AFjQWoSOVBugsdQOAgTuTMawIyDxaVcECfQ+J8
OgVfT+Oru7DX5XfioUxctoJ9nmoQaQoByugrqNCloiQ91E0d9jM3FGpfA2E3Elh3nJwfNg7WnvLs
XngWKIliazMzDucJr1LVUprUCDgcNAMdzPzdnKz8am1Oj/pX++D5ToqezS2WkGnzOQHPFLuSGtB3
fC7ATHj7wDGUZZYbkMBJ8ZwquHzsG+ttCGMKthXtumU4YiTZOvTnUH2MD/i/wFTIwWqHtMmtLJrL
8SM4T/qEUyu9rXOJuHLf/o7PYxaL583Y7xVKrBkKtNrs7xTdMUHjBBD8WSodg4ykPSg+pKpWLygQ
qn87nF4E79+O3O7qh/YmxQ40P1QU/y0sHXXPDpFdPvHNGOJj6GBDgDHnM5+TOmTI+b4ft9nIinFp
uyBtbVyPk/l5jm4UZ9zkEjNCvTAFHj/yysaMWGNNqcde87C6hk2HS+C0f7HouGbj3h+vi11I7Xgh
uHqUCzv/bLyrt5dkA4rvVam9irzECl7plXdsnMPgboYS5Nw10Lfq3ZY0C33LTnLu/XY2jjPjVq63
SUEd5KNlK1/Dy6NG+2BrqKXad9HxxYnrG5EFhmXLm1ZUexUvHAKLcqdJxV0TJsYvMzxljwYvhzBO
Jb5hMiSNqasvG+QcUeZJygOGKrSNszkvhyH1f3rw3gd0s1nWdk8iD0F4BqjRLDZb5WOFqXg8UM3a
V9k4+8TNGx17runDVo5jZ6rvE1ExDrhULb7B9ELXillBMEkSuz+6aWlzXSoO4wJqtCl/dOkH+J/M
iMWuScJkPs+1ExZ7cr2LnWyxihfYF29nwpmpBBI8XaNu12xbIlOmIgtCstELjIFfcHy+1k4oHgYW
LsJhBzn42NxHqPBgI3eDh0r0M/MVREbyxBCsg4LVSiTl0JOHFWlTqpQ1cNFR0H9axRmIg3a1ZzDA
AFrmgFSyILLXY1eeRr4jLxEUzY5Q6svxQs+baarXjgGZ7uLGpiruNcKsLQN+qTJhaY+s16iP/MPW
QkqoJgqGvX25Yyq6sWxe7EpqmaKgNM/k8q8fpNHm6aKIAS86N17qve0el0mRN3nhzr5gtdgzJJjg
Y0JXl+kiF+N+CioHu0F7lGB5yTjcLsERjmqZByPV2V8e5kxrRhqdriZqN1elTOU6hPQnqF8BlpaG
VEv2RS5NgR4MRRABxWVF+1BNUydiT9zkc1VAWB/6BUiOL6WYREix6xMq9WtPD2ljBZv4iFCCQKWk
XR0p2OUIHERp59xhf8iid8aZpiBeUPACgaowpdTRgrzZ7eX3SzajpotIwtcDMr52bIInsLFXhYgn
X+eRbXZe8XGt/ZQbknhnp5m1GTn393RbXdMes9jxn39KVmL11rjy/8qhz1TtZ5AJz9Zfml1rWQiC
tTCWGsVD6iE0gMLag8GjCsgbjykdHcvOvwU51TbVWfwjODD39tl1gyZ9WwGlxw1zEVFyC4aqVwHJ
93uVJTbFDqUVXlMfn+c/rDHdhVysTPLGs+3CcTV9RIoTiMkAMX6R8ROZMw+48yMYxKjVWEpqM3l8
wwgPbS0i3SlCd9PrzPbjkv6O+FUC7ZM16a34tFEvPYPf+RjZXkonp6nkxP4L4vO3twc9UcXjiNo7
cBmYMJRvPZr9uU3ESbLFz4+jfAbnT8wCNOKou3Z4L9C0cC7F5Hqykkew5xHrJX1yLevhT+32fCrV
Xz8xeq87uwyC8nQKXEajl4AIV6BWyzswTt4Ky0H6jVX21pVINHAoiISegFKmwyah5cFvzI8d1pJs
wD/0d2mHkpPOhzmAxia9sSD75soO1sPcbblad+oX3Q0uaLB5l1LKx3UsLJni075j31CARRZxmEBA
oG+KbL8LaaE+2giWXNmHzDE2t0ZVdSkHNewLCRpZLZ42bxSr3lZnYMRpYDzu3jQXGhmtmuwAky3W
Tv5w0OrTdn7B2wv6SQX6150vUHhkGPjSbfgWHG4q765T2mJG/yJSJic9yENOPs7RBtpZRTtzc0cc
IxyXGbPnPswVJUl/sPmY5l5R7DBRwOYvSlE7PM+9s2cuJn4LyEXVwqeyyGuGWqrMEZx5eyqCXm8I
op55Dt7M3oOIDjYYeTbjbDwsHc17i6QiGgiD8Sg/Yd1RloDsjTkg39JqbypjVs3ABvX29pjIvC6D
bxNC3IlfrvT20/CNjlGpiy5Ty9dJ83bHX9ZA0TNyL8mRS6nm8MO8vcgsE0/36EihrNW2uzjrhPn/
HWV7CSOL1SyxDmgfkDIGKaXKgGK47d5IjoZMwxb5EeJqq/i1ji4AksHPQbRnXIiY4RDIItVE9CIK
RjxJ5ay66rKFgSmrtE1y6r88+CMEF4QAKKpFH6+DGfhG1iUIa7mVmJwm84pijrK8p7MtOr/kXNGw
GaUVlwIi2Ho/cQbN95oqIFqwXnLR202D3YGwjnE5ACD2tdcKgFVWBDfJDWdXxCSmdI6CUoZcRQ3V
Ro30Nq/lW5lvzhjXgDRf4/KraTyuG+Newv68oWQhN/Yy7B5e9XwHsWnT0wUZuvVuwLEFJD5rW3wm
Yy8VFWpe/FslO9KhhKqZpGAYC76NUfBh0JfHpHPIxv3+sT5rZiHQckA3HmSqiCU7azm2bHEYZER2
/Qqf58Ze2WL+g5qdc4NgMiuzgyDJofU+AfOcVrwm5qJNxzjZzA9uzuj8Ql99pPXLS/IbGBA3mP3v
0ukzGgiZgUz9aKttQ+jiL3M9+0TVSka+i2w342x9kvJuwAWP4xfTfShbWoD1x1/86qOLOozHXU6q
bsg08WkbvDC4P3s7I9An4MWfKa5WwAsjgWQTyaKZRvBmgGxq3Vumv3nFTXdzietNDZJzGVzD/upk
Cq3pIdoO0eP4FSb9D9jYWsHjaQq8zw84ljZAQezNvB34GVmjhuDCtwgEvGrGMO8WSVp8MXSrxo3J
YZz1XamzDZ4Sh7edQcMZ+hnrwvD5bhcYESM86ORSSRs6WqZdrvg2bKLIqSRFpjyU7lRI/gH80Gab
eRiUVc+XzgczN3DMnnIFVHHrkhhTJQ5pUp/j7po3abPXJnjGChNxIkOxSYQJCRu95RPFzifEvhsI
1VUJTId9L1zEXQUm4HTfXeGN64K+FLaHmcO7/e727wWJ1lIICiWRe2u8za9NqOzjZBZudYB/ib/9
ctzUnq8ijrwAzIJEx61qPVzf43PppmQ7MSwLim5x4Nhp88fsOEXQOLbH6vRToyn0g00Ac8YQ5PJW
fD2un21h7Hsyyu6ebaGqlSyFB0N/DhlExpsFvOFDSC85542yJhp+4LUXHyMasY3MGWdbsciiNPFX
wWn2KcJEHFgWcKJv2lg8+Twww4rkin0Qb737Ag1To3FlRTaTRZXoFhoXMV0hNQWxPlTE8apmArjY
vSWryKrxVGEEBuBT4f+e6yZMZwUIeEGvNHmpyW+ucSg/qCMzr26jXD8+6kfibC8zD1yS2+b30HhX
W+PH8UWoJiu3YGXXl16MrslKUbLcUnSOGXoD47Gqh3uphhdW7fp+nctfKMc1JFZI5n0fqGVJfdmL
XIJiB1Jl0itElzcz7O+QooZb5C9gar36kGBRUlHmuBLI1CXEtCeqo8ohpWdm1YwA890k2q4tZcCe
jyNXjxFagp25HLtrPxAcEXKjXnsA+/s2odrm3rEEtDUU5KOaH4PswW/0YOJw69l3dA0hagkDXkGX
v7VB+5iwNPHJIF3GQHqkUNI5wdntUAAuPJise5kY4qS2UUS+ImAgNx9Y76b1oepqPX/lBtZjtPRb
QS3X9E2+2+zKKasy7TO/OktYD0czkFmnWQ1ZYkaxVOtX4B/h4RgwT2kl9W48JrrIFCTp3Jhl+K6R
tkUpOxASTZxnH8a0d/sY1c5Wjn+1FEjWdMe6ljZB6k9QUtwVGVTDGBsBgjhg3+tDku/ttP/t2JzF
PxCCiRGxo7pgQbRxjfpdIz/VAiUh/ENSMqYRlsIKw9AHoiaWMgUheKZtXRu6WF/cG+Z0ZIcMtJnO
kqF1ychMZxPzEZnV13iEcFpG7ZkQPnbPhsUmHCWk0y9Vdubu7wyljbHILOSgJRmmuFa82thTQ7J/
Z4w9eCioF/F4OyRGer2dwOOgu6vnZD8wnqfMDRoNrc7nd0dvXwcC0fLTDMqtZA66KD3OllNcWup2
r6dMsCFbASqafti8WY55u/4bHqNH5bypo8NjaPpxxoewdSFCKHu01aOcRWe3lzfhrVIv7QUMq0EU
iVyoi3raCWwKeZm4Nhi5zB7nZP0FJuHoYGwbRTv9lg3b72Z9vGTY5Rc2ORMAf2jcG/JdqxmCU6YB
eluaVcHxxGrmmkvgIG2jt3OHt9rag2I8l1ra36QmAXgr5JZKEHYuEmb70AVo4+XetGAkoYCcmvl3
F2vFeBsjBrLayjyYdxKZ6CIWezEd8A+FXzvAxHzh5mNhw84Ee6r0M+9ihvW3FuT4FuFFpKf4dlHB
HkuUNcaZcyuh/VtiObiqNkotrp8eVNKT8XtOrec2j9ce4L5ZkXXOQYmphxQ1XZEXKrjBNeo5knQ4
aU+AcBI/CDAcsVrxp27jG2yqhNn2+bLmKt7jWnBcX6PEfuDUqMdHNiDcDIwYGGQEb2mZObwlNP3z
+NfgoI9lFZiOU3oRoPiX3IhadEDmXEnQ1OBrISnOXtKWl6m/icPvT6obKbjljd2jtRc5UFsDPNls
jNCeQu5hIF6YUA2QgPf6FhryDHgAtHtsSlRclppT6ifXfkMlvIffhyaLV/IVDLlG6i72RzEaXLUg
dvTHMLcTTuAlsH+XwEusxYow4FiRSOlpL6dKgwF8LuB3/MZjHxgzvJ6yLeKhrzQgg3yLT4HtbAT9
2pbisBo0E52IDc3sOWLMueUx1CoAJNrVfl6HTOIMVGQiqU4JNJXMF1XL+4h7xPYW5tv5cyRrGqu6
Xtz7tKKT47iP9xXTvsvV85p77OCmuJgwebREdNgtdBM9rI0ydADpBN5y7sB5d5eWLVebOrPhCrm6
DNZDbf+y6LeyArCzEKZbR+/fg+Bq7QUKvaIvVvL324PtTCfdXi3tYeNpIvmmkueH/g6sraH27vxq
Z1rLvZXqRwyOxisbKFcH7bN6yB223faI4FHL7hausE5AV9aEAGp/E+j/xw6HnQRVqdnkZv4VbMX8
VPtH7q9SWljpBnA9ObGXIqhQ+wR2uZpBSJrSTi8RZDYrDiu51j06uj8/ZPQHc5InkhXJg1CuWGVr
qYolTKkLS1GxzzTEPiFceja7w2b7VTFm3Q1RGV+LOz+SGD4ow4Pw/e73EQsAW5o9si3w82QxUJk8
0pFHdcKDhF6Te26Xthn0CO428GCOBYoheHqaOZiBjUcfFyn2tUo/rjYyuCFter6CdnX0CaISndzI
kQqodEADr7sqKT3cgBLgi1XkaOreiGJyXKktTfWLRQ7ufE6QN3euBrjMdWvjbmFIHJBqse+tbwbY
pS7H/3SmbSwT5MEdFwHrJd2VRrD6XgeeOt1pWn4rqKTMsKCkF0tA6YYqFiTCY2SF7SuSE62Od973
3GPwZrUhVbikDeECtF8g4hZKUoeoiwTJGCfctHfJ+hFFMSE6jL+/udNsDJbZTiH8JrqiAqMZgfpM
emBGe8iB+0wEWq0MjYSk5z6d29BjJFRBawOp0mE/N31A3Eq9EzNvWyF8/Wt976oFSpb9+boNJggO
eZAzQmuXwlwtN1qrMCoJC5KLZlUMk3ZV1WwiLv25oDsaQQLzQBULrYd9hzPLClYyi6DUqKk049aN
ZgoaqHUWkWropxf2hAJUKRRzyWIx+4nEP4Mww2ZN4SzSYWpcr8jg6Qo7lpClT9c1qevQmXhQ/EAz
UqbT+84c9aEYf4OKWQOtshAAoKewewp64UNEL7W5AFNeLIUs13dvzxgINV68Pr1v25ls4B+FFWZF
yGbuFrGLzCcGwR+kz7SMCLJaXJKPas3WRpUwRB0KiIKKpT39VEpPZm4ITF18fds0GVhGAO1L+1xz
sB9pZ1c27vfrAxEeQN850kLiULT1kYUiF8ALscaPjVxJmAd0EhOndkHus1duGYjetmVx8sTdoIgu
M5sGfslb3HAIQif4tP6qfSpK5jsH1/9zoGn9v8r1vIXV3jYTsm1nzq0ZBN61GAl2g/POyHD/9/yw
S67jnhCejfIBBWjPeC+OKlO26c2k5zbfFjsa9tfeY+W+5RNJ4xpDUfZVTeFRLmbTygUqMoYOMfqw
fY86couQUtkrTjLIveZU1NZKUGWZg1kObh30TTDlyM8brU/cHcs/4xQFicPGZ2Aq13OqCjxm9I5x
6yVwueVWaNB4W7DmdpxMJ4FSy4efKy3gYiaeP+xB91kj477dgpa4TMzESkhJE5yqhTggcYigLHDR
oRkmE/rvn/ELJyZSFO4KbCuow2Mlc2Y0hN2RZmpiFywgmRuzqRddW8wtEEs0rq6CryZS9ZOmUiap
RPj3e6YeZB+r55pmh2mJ3BsbbqsiDSHhnQFLRs9NL5y7TI3jHbNAiyL3LLWXZTSKMsoTUu+OVeCA
mj1xu9vmI7eM3SmWj5+/c/P+ZI17eAMh31Xu1HYkQ7qv1+HzrUz99ZEdFDs5uSHAkNp81Qs40ITc
pWPiP+460Q+LeyAhZpWWxsejoWORtjDP6DqmG2CnmkqAzskGz+cI6aSb1bB9m39yiZ6Y5CDLLUHe
jCt6B8AquGpUHlN83Dk+5dhZxMvlFr4DdU/i2i1QC7EihSk+/pA3p4PPU8jr86q3b1P4sFimHZmI
BF5r2CtU3PL9butWEVCTv6XAzb+KBIXQpbEJ0/EyKTgLb+U440KobEYnZo1PbTh0rBY4LjfpaUlM
C692hn8c8OulQftJk57jHmYCvPYmcjnOW9oboPjRDfqieHVndv50Ev4jEMcaQ6wPs7m7SxXNnH5M
FaopmbQa97wTwduFPa3sa6L+XcCQnPH+Hsiu4jrwncLfajTZaAdSdQZLVTz7WmI1A72smhJm5eGj
/0D2BrhvHA8aGY/n/T9/eqY626uA7NC4dBqZQ89eRdAX4/SGAeB6dNZbbztfyUW7xRLoIEdn2hb4
rbUUXCnKjK2pNLsotSuGA6swCqu5dFXEi/VLFbh7fQn1+iahUr4nSqqh9SigW0dl99rR8qmpgVA2
lDyHOdiH7UP4kl9Gesr1dLM/+yDt4C3VdO/Rcd+F/ytiGw7PyzNQv8an6AsUDpSF6CfsfdeCb7Gi
7ulBKpYxDPhzMFMV8h57pAAxnc4rFqNd0aekrgrgA/P/q5NKW6RVe32AQDqQ1NR64HEEL+0oKDTx
pokPcJYs5XVP3npwX+4+/D5K+eiwPR+PKCcEVZeDuf4dQa1WZiQ0U5i1aSj9XlM2tf0t45ZW9MKI
dY/NDs03wwjLg8dTpR/V6UBE1ulpLqsD3rUs9pLXeNVpXpU5yQIm0cURx0a9GhMANp22thaN9ngS
NaZS3pt94w3sBodHFKh3/mL6W+JalfA7IJ/oA0mpoC4pZ+GsDZnsi7It5zlLLVC270QETCaz2qay
B3q4IGrFX7aPMkBzmxuFFgPkKzdfV2/Q51oenMr4RcGcigRh5LnRQzPgbtrEDnyIlYb5qyBjVQAQ
hvonoktwaO6I/9WN9lqO6ItTPlw1n6rvq76otbv4ASDld1VoQbb/LY3k3h+Wph7KwTGR4MYqVa+z
VbxBgGrSgFyDzPK9YVpb8Wqmb5CB6l9TH6fABhgTPLOEZKnkLAKdsMlh3qvorC36Ha/Mlqauzpcr
B7mbAfmCe4Cz52xeQOxJr/vMeVydFQpIy/th2NDCiwOVO8ggF7jb8UL9LAxH4iH+AHW3Qfjr4jQV
1YIR3ss2YSsQaQYJAdl9H155gRTMx2SgUMPmLpH26xdH2lWeWHlSySwhM9+KgQbUVtGXmMeM4rmN
biuS9DzvQi9+8U7XwnBCTbOqwZjr16GnqbjsL/4jkVsDbWFKsv8MMe8xYERxQ6qgV6x6zjWa/87u
Lyso3bekG669uOfOyu06diCW2Rvhi2pAoJahhi5PpZ/8+6r5SHIJblOMEMSw4eV/igET3SOoASIh
vWutlRy/5Y4o4+s/aWeKPe+bhjtzSK38lxZKSL8o8mOXDDEdBy0yTSmWcYEDQIVvxGMY8O8GTaKZ
R5mGNt7TLRSopHEj75A5LPIZPEx2e6QsupANgTby3z26p2bkKKf9xsOmCR8bs3RPun+kZ55eq2Xw
ni2Nu/8/guet5UUpfFM/B+c3dj7Q0SZad+w9iY9NkTbUVRgfmHvNw7Ye4MD21gZUIus/EUdY2TAz
ni4s6RQn9CpvDUZKjTMQfAUWS3fUAkum8V1lWQuvmSXprQX4L6Wez1eaeRk0pc4xb/+7B4PBkEPI
Qiq4nUgfDvQ3ZIhu+Iwt8cN8HjbgYKfTTP477q2TN6f8cl78YFGoKBOeld7Y2y7EmF1aOUshZ5Gn
+Lj3fGGA14caPFcw7XXUm1u7tBu9whftvNDqDy1zggF+aPXaz0fuvdGElbEhQTtlHXhb4eu0YJ7N
xmK6KVzeoZhltUKQJ87IQibZPLyvymLsJMgYVgPqptGF9E+DCrZuGZtIKbMi6MNpc3bFisDS9KNS
6+APxsqGQXBNaM63z1z7bdBRgwb9d92RtcDaX3FVON6WyPokQefNe6gijsTpogsHA4lVZDFmOt1y
rUwK97nCSojy6H74epFsY9a94CZ7WqVNOUmBSlf41wH8phb4KS1D3yxQJLp2duqhzeeEiCwPLMkO
apKFZOs0YwMI+kcJCKq0PiONvohyP1e/H3t3WnB71zzW5OXVCaGWJ2zYRnK5Vrl5m9x+Ycu3L+Do
xrNwj3RMcqsvlxQ1fxSKuaT3aAe7d4KIV4y7c8zUfe2zXCQhLKo5abJzrp0rU78SD6TFIomyNTMM
zhHLrQcwMG2LeHOW5k7e/TlRpNL3FcnsMZFnQu3r2EFx/H35toPjrEm/xWsvzyyB+O23nshuVmpP
U5xeuJnPsCK4ULedoJHGivNBM8356Y5Y+HtP76GI+O1PzzPev+gCGt9Lgz0/A2rhp8V3jGSl/TbZ
JhYQNJCQ9Xpbc4s5FtxgGNwzhpvRYJdFKdFiFkHQE9f6ibLvOu9YcOLpMcKSqwxZTz04BEpJuDf8
OI5w+2218hzOjdDh9HphWVDHcRHQZs+DL7yEKclXu7njwG3n1iMFS/Dp5DO6DUoSTEj+dSTZuD0f
QZRhc64A+djYnL3hB5tdzfsqQ2tsirOe5uWWpKDqIfqu3obErzjdCCaxEWr5t+MihviPsWqs+Kdy
39q7ko54IgHWW4okJOrRm6+JApQEqmhiZIy71M81/cunFXZxMCK0MLq21cBZD6byJ6IDajuSEeDY
Ft1WRx4CauG5qdUlOzTGnyoFwAxZmA8+49Ia6MFLjBUs9L6/t5jrrXYjohY/2EmwfTjqxje/1BT/
uXgDI92iXKe78qQXsNzlaeRvCFhwzcR81Okvn58b7CYbi92BTs5hPMC+YFRjqIzmLhJDvdUkESKM
NEUz1kwFIa9RGQjedTinqJ3FdaAELkRQzIJIbseTyRTybxfiTdJzcxW+77aX8icW0DffCFPY9oPR
g3Ka9A5Sc68T45t6d7MazqyOnb4ZYf7+I+pwWqZPCqRh6sT2j5DSAzyDaDzU1MOejTtQ+v1Ydzfd
gFULfGWUWeYZp5X+u16lK181OGD0nN9DMGwXwXxzcqAPw9qkg8Li6GvbDC0ETtPSvIYs+pFV1so0
/qV5GtytzGlCz8ypRPH+CNRTcJydzCW7+mxiRUfd/gYP4PrcTydRXgj2N31xXvdbz25rPh/vNbQ8
NNvZjAFACc0LsgfFTQhXQ8FROtHZKHXWwx6ubdPs27cAnV64EAggXL/QUXny8ocoEP7VxyJArsMx
wZ+wF5nzYdG6xFWDZNYuHp3DuJbVVKqr6q+k13mFfu5LDs0PnNOGhl4yaP9Ccvb0mOCBzz8B8Vou
OPNkNA61kUPVvf3mzQcNe8xbkFjEQGH6QWmeTCNdaPr826wCstuJJE2Sa2/GB9kbD6FA3riKV4wQ
s+9X2/mgTTU6UQuhkXZYojUC4s9MDMxiCESUCr7BvGzrF23ySnLCP0cN2ADz8nUsObndWk2kxDE3
8dI4Vm7HG9UpqzbLHwlAAc3bFLXOAuMEoCh05bhfUEm7Qgb3zc8p0uEliIAfM2m+UbPPSZA6MYd4
6jXzBvjqgmvlGYw81kHE+pb5aeOoEVAOX/NpUVt5lvkdYEPMdsXhtf9u1pH7YKbfrDctdW1AGHh/
FwAOzPKAi/7xZYGqiTITKkP9t59sSDXAk2Fxs6ZiXWE6R/alikn8EVfzslWpAO3VFRtYqOkkodyk
17xwZoyfjBJWEpRWC5nbCzTZfNJjWUCZ+lpbfXFNMjbFXgBVFK/ffHDoeldgFdDoHAx0wcTzLi1w
8S6jV95UoaIP/8pjB7QQEB2m4p7akzcMkF2aRy2CvrGtyb9IXycs+AWHvMHz2nWCyP9FkVNxfsPY
chx366AkW0oL7M0KUr3oY3IH6NUdR3yF/0SWCyexKPCTVQHu6k2gGGXlT9aPPCO/+m/Nn+ju24Ws
1vDk09MKFla7J9XvUPoR3wB12Qk0VLM45PazIsParDABjOxlppCphtZ5KjemJtZYz1qbacap1o4t
YVxZX7xw00i513p9cXPa6Fr632OFW/vnJuInllPf2x2XiKA5awvFjpg6Qyzir23Bz4bKQXGhIrZF
dqa1PT8/K1pl+rIqEn0tqLjL1at2qfmy0DUMsXU7isd0Luw0Y7qULWKt7qyIPX+vzZ1qAEEbnqh7
CHpdV+MZRYQqUI4ZofhmzZdWIc9VOJy+s/dlbQO4CIEQvbP7d+0XTrYxzDxWET6DbFED7LnSLBJ8
WTxLX1aaDRIEN+s7if0U++2HOtdbg0rzLEm7TNWF/fpEfVi1oKycEFeFagJ3PuiQU7Q5p8SZ9HKw
cw4UEao3QcYFhAQrEkEUYBO70vrtQpz9tFttnQGjNlolzu3OxJsHUCgVVEUnUVR7GSC2YIeN0v+f
SUHGquvyK2Ttv0RdFybaGihxKORRB1YKUltE3r+YScD1TCgMErIWe9L3Rcrs3lG+9Lk/EKyQcaJs
Ew6fzRB/ffSG+mugm/VKYq8mokNjN49Ej/NncvHK2NGo5g5XULWEyRBmCcNoYzsx1QHDeN6YKUFl
IdQsf5H63rvMmgmiDAKaVdw/+M7HgRWyD4kg7LvyG70mpdjOmEOLzeC7bPG5/ZucwAtSzk8PShVc
eoUAg01qxNLd+FZDc/a3Q1gS3V7HVVs97tHWLf56NDM1i2XEzNn0/9+++qOHgG1gjIpiVlgJNndR
QGqbfoM1jyq/ODkehnRZnebBpvPzWUisBbrLeetpI/h2qSNocJGsBir9JzVa8NqsedHdaDLpQrqI
AjXLbBXhWq57DFv96X6nTxUcyU7wijym0eZmzXVhvrQGQ7J4zOk7YzPTcyvoZluYhXZ7uUaS8ZPo
6e+yegHsthQonPPsl56C+2LVw1OjwhVurtVuBL0XuOm7e/Gl2Yc46XJaGmEAjVlipcMy7W5A84qH
pSYXGfyPVowUwTvfIGtuyn/RZDvyHscFRnI/ZpGmgGDNAUA1ziqLPWolyNUDd4NDyl9UiyoaQWru
JxTKCXnPWzfaO7O9Fn1zLOfCilhvHrHSTrydyvQZmf+o/7Wp/XrKVVvEdiAaHEKwvQYlQdLEUHgQ
e2WIp4AWTEgid5Cwbh3GUt9OsjJYAXv62U7dJULFACJJZL63NYnzNngP/y1f+VdMca9EYD30LxMK
CdWUaW3bdyDO1kxK7hc/Lit9oExz2CbFvOr/JG6kLH8fv7yn4updFDQxwhLkLhmsv9060AmC2vN1
90CfTcbYvDNX9c8wMF82EZxvdpVpFCjn1qxelbtgTp68U/Fk2bZ/Qmmsljkw2ijIKoNbJmNnukb2
ZyWC1qRCnxFS0tsBs3LVqCwRkPgOL7+Brb1PXpo4DybMicvY8RzE9U2VHd5jas/4OaZC84JVdvJX
gHzA4+LsGgflnCvyV3T5CHaYxBjO843kUTJQBZsrwUSs6NHiTiR53z5FNsX9amOivtbSDDrmXH/X
4djaMbmFzs/OObiER1TOhfwyYkRsrfU1FiwKKV8fVGMdY6IWa3Ht1bY8TGetl/rSmqckIKYC4b9A
xs/VwPey2LeEWr6q821x9d4PVrZCslqb7QcT++RlgqZ2Kb/iQ2sZwdNEU38C5sV/PjKSL6W7MQN9
iFu8Nort27GC5wsQVZhRyNXCbDV+7eqj/Zlq063m1cM5aAN7l1sftyFTyU0GBSHfCA5cSiuQDMsv
WMSP+ylzGqWvNq0wpD8bxAeBbJUEnLEg9PF6ktLP52S8HC84dfakCjIwA3WkDuZ7ZQgsAbEpg/A2
9SvuSy9xJOhmWpBaqCEsTmHMs1Dzv1qGEKwFNLLvPiRS3zA82+y1LubiaC9H9MbdYduqjBFeCFEa
IHjMQrGPut1AJVcrhVxKukPHOcYfl627KcDTEdjtIHGJr4+RG/+xs4N+cQWpYy878mx+k7K8kToA
/bv/Hd12/31jNBDhJta6TxUPCLfx6d8xeBObjdB804696BZ1Qlzit43uWzoXeq3VZVGFFj09n6Td
UIVyX3fWwqsddpZsa1ZuTjr06gb1F6t53Iqg5VLsohXnMM7FOBEcipdiUYzQn++n9FU8ho0iXhiv
3tc8BD+3YqPWlxvtD73npxVSHHp2ni+bCA0IgiuCCx/WEMM/mrHuAgoJDaRhgN+4cFybUvOsfkb/
6zzBGbLRLOugKNH6Ooz0zs0j/8OYGrmSxlFLjU9NNt/gIpuvF9m1ys5OalpRdYZxw7xTRTTsbj8t
uDE0t48k23knewdh7L7q1tci4o+1X5Iy4+O97ZL8XbpJcuJqCYcvs8jnKt0EvkMlZk6g/rtPvr9v
EQXqTEbafNBYG8LM6v5uZYS4xjXtCtg2zTwmWiuloMZoHNzzy4Gcfte6uWkFMsge+ZSMBotNZETB
wBqiVg9yzSars9igfH/Q3G20a5FPTpecPQa5cbypqiz7Egqg7DCjZmgije2yntZytKgjKmDObR+1
wPk1IlGQ1B/R/PiDVxFn+QBG6zs9MneBA/NBjT2vWHhFAupVjZqZooUHwEz+73buI/ZpL7Ag/N2L
A+AGUcRscdF0JQICmgw6W9BuUbYQ0BCvcbVfrc9F4fX6C9dNxmIcI60dXcqKN97yEwgT82VwSIAE
htDhkjHCFcasM5LBbgOu0bEchxLrdsLUo02W5+qA+iLq+By6gL0AOXgBjaVOntJieeLrADBsy/8d
qTbHQQxIEVQ8WukxrlxqHN3pADaZu1i04Qy6Q390PaU+VJ1uZ+efkJ3efkIEu14MPkXfrMq9WQru
azsBfP3UXZH1mtPfQkLMud7vHqWBHbQDeH+RKUySJx60o7oMQoSJJ+JvRE5zd9U7JkSI27KN0MVW
T+IA1trSVSb3x3Bisq1LvxJglY4ftInnItYqdICZSutrRGJ/7qGB6PSRXTLdqwEg4s75op4RTw3k
MNYZNScp7j62RK+sV3lHRNkzTO6J0VapLT6O4nbDN+b/sQBOjbtKitomx1Qz8koxkLANx+k6SooP
9gkfGcbjQmgPzXU7WdcrRpZHWgmtsNJM1Ev30Jy3jSCnIW9WHWzyBy+972c0npWbrGLRz75MRtI5
J6ZyEZ75I9ygQVxKxB70xucfhlLh47+tEbisBbAubPzYhXb0ZTazDzZQLAyLXe9ABEFgNO41h3AG
FtgklDqnl8BdiexFcg+6sQbsRWJ+ljyP244NQPp47TydWAOcTpbo2uI+2umSr9kU0d6VQv9jQ22R
+L47ckyS9whz90851J582IQWVQFdb/tV4y15J/BAIIP1EjRPAmp3tXlVndGMMnZ0zbA4h6JKpXCA
F+XrX4Ku8NoobbhnoAgWOFsYoQT8lQgMxAdj4jmvMiMW/2v/7DiOIYwpZE5iK0TP2K1NZeJIf+mB
QPEAYyjCnnTH1YpROPqOyg/a/kDPrAvyU+5qu5HOpAGSEbbteufwn6KqnSg2YSiQaCMNfn/SQ9kk
eQxZmI1Y57mKLRo7gzflL9sxLlRKUOVSzZ1maBnnz7OVJdkMmRUp/ZAmb1h/AKeVnBuc6yg+Yn6M
b4miRJucv54J8xCPxgPbv4qMkZn4Ztv3NQlgPyyM/lvCOwGZUNQAZRalng0MEBTgoAXXLoC+Fx57
zB72uLm0YKGYZVM77KQURhl3+zLrY0XICA1v6MMjkI09THznxalZQ6JpbXJ9Qd8uzIsyItBQDRr2
So4FiV3xvrRj33OkrdFxlKhRe2fB10FYWfTJNAYc1idpDoxtLel23KtfhCqyRu4ai5BEJ2qbcaM+
hmOqyN4jGvRIILJD46PWY8HTgRoNiKv2Kzzp9bwQWSkQkrkopJLV3D8M6CmmgTSvYxg2ucUv8HxR
KZsqi6nnndcHpGnnY2KxPfao92K/atYk4UVbQmIVhO0C0eEAoIfltBZZ8QBN2e/u+OwdcKFq2kfL
YdrXIZDvsOx23496EjSKGGVW5IpPrhfJvCr0CtdSGjkje1ZgB4opM2bBsXWaraUdXI1dewS2yi8a
boHq5hhvp2BST1US2Kj4Ey6CBUKKXqq7DB9BzQSmobJBjx9Ji4lsBagdc9ZKwMIxp12kjQ+VdSR5
1uEhzdNKIKOC5a2Z96fgNFx7tDMW42qNYNGJ8fluo5JPqTLZrlw6aJzWZYzN0p3eVdl49bAyGpDG
B7YVxVXBU5HpU3Tex4FN0dFf1oDWOcllv0z6iUUDuaE4SNlBUUHGOTCLLKHolyq948WZugu4h/yu
yKbeLKjdaH5HaOcZsQA6pCj19qdJd6pykUrL/1DeH7f77Qllc+bLwQL8FrS8qWc3O7X/329FlfaS
58p6RtpN2bMDZdXFwWEH1MHhC/Z5tzYyPmdifoiLyub0DEUe0qoTuORVsVxU9XY31NZB3NN683wM
Hg2oe8hgfCEtIjk2Nd19z70YGKcU7ky+VnMSdrrA6zYMZlfLzmWiRpkkWpGnMGSiGd6foDIcC5i9
BZgkTbgXg1yuu5pM3Y5Klcm0zzCl6F97VpGvtoVdeulVUCSv6HFdLJOzyFoIlb92J0uI8oc7ePm7
a1A0cy/1zTlgAfm177m4ERQ4E+bxVEt0U0Bf1c34TD9pC/rhhAcaP9DyDtyT2zyagbxX9fS8vlue
JGitnNG3bMUwf2XJ8o+FCPd0BbqqMu1WNhXAxW4TCCMDYbZsGJWvqAFYMZI0ua04BJRo75f0O1tP
CuOT+ADzJ3JH/JZOJ1K0jW+Mj70LGUB28CbO/tG+naCIqwJoeeOkvBWynwwRbWRlpS2+XtxIVtYL
RcupAyHZSMHOnifjp+uvqcuxr37tBp0WGaj0ufmuiX6afqXfc8Dm/7qVOkBUDbX9U9zvJRBbGLz8
Dn0bDOed9jcgUsY3SP7xpzI9OKzaH8qoJpPiN3r4wGezjEsGbeNSKmtmThLOdkQReaAFsZ9MT+Uh
syzv9GPicpmMH4bgNYednfnB22xiP7UqVPF5nsSq8siP0MF/V3EFpRgUFe87s6jMPdsRzZXG3TDJ
lWjQHsQ7H82S+sVe2erqlvfwLMrhT/+7ACC+w92Q9m0D9Z1qJ0vJecXeMtp5hxFt9IhM9cwlIWi+
IU0mkk9yIH1VRw6Gn5jOzj6XFWR07AHJPh2rRREUXa/5wcTZC4G9pGzI+T8TycqExPfJmQFdHhUS
qoGKGtwmDv3k7XXISHHZMys1PJdjk6//8cjpq4y9pCHNsShozK1rCgJQaqM4pHZvCAAaAD7t+Sff
61haFl4UMqCKvFz7ywtJvMvX7rpwYN6G4nZEjErFTi+R2Zzca/6f8X2BxfYyAAAgjbYAtN2LaUyu
BDsMnj033kVDhBv4KEhZS/YfaJ4sAjV0zXN2MOZCzlq+wQp2+MzKgbO33U6A+V3SVo6qSwD2rtTJ
DiHUt+U1KWlAVwm5S8fCtomHgd4wqi5011/Mkc8YBY2ZSfcaqa/IGDzsdZ9dnXW97rTNJ0KDYIg0
cll66YKiQVjEyDJQjg1A170gUPj+FTeuZSFHQrDMNpngfu/lpjmzZBnkPCf+aW4cgZbvU1diE1fX
rMvu5sDm8P0cX4MDY7hQdjvBn1Zd9o0Nd3Hl8Nl6ub7PYMUKlTIHSLZtjTfizOrmr9lZOR/VGxk9
NK9Uli5D3IKDCAGcC8bo2KZV0z5s4+ZBptis7lq7axNs/c9FeQjxeiTdAl7VHyAUn6s0lAgTNzzL
nhIeQ0kEDq9Hp8hbHSx81agsm3VZdAQQMuoRzSMjSJ7anpq+EwBwov3kM0VXnXZmcYNtV/EtRP3A
mfaitH5Fpc8CjvgZI10GcAyVNpQG+WgGryOrYudCW/VeTcC6WXqJSyw4sAb+yNou0CNM4Gn4vzkm
mHJ12vKUytYjEWhsGQFIYK8hbHwLaNMKoyPXaMJCxjF4mu6ksWn8Q9DGntx55+Rnb3toykwnEIFr
Jc7o+WdKit32CCizgVJs/2Nap4MS9+0YDUpu23gcHNzQJbCeGW/WfMvpQn23bnqoBrlg6xGBj/x1
Sx6sh5NpK7l+GR+LS8O25iejzc+LM4ySwce6heMlxzKVVdPSYawFq1U/iwAZG0yOKqsp1x5Cr+sG
Bup+8AotShuTTlLy6GftsQQGPNd9dWYIQY4tgVXfj5UtEEDMxWOjHx7KGiqXuR2rYVQgwdGyROEf
MwZTyXFoPMq0t+yetSkGtr33EmnYRhWHlNKPy0LokL+a7ci34vyiK3yNLZ5eJx0k15MKIdetvFP/
beTE5o067kAoJjirmXp5qe9/ONjxeDfomgljaCfHg4ZRG4GT6PRNXwQJlw7cGnYPu63ChybR7yHg
CudHOpki3kBbnfu122E6je1Y/SHI0mtCnQ1/vtBsxpClkNikIvwdBAIUyLSLSzDZNSKt01TSZGoS
bxI1nXRe8nb4XtEX9Z70SB+6ejyEOn0osGMtl9YoOXL3t8qVD3DXO1ZfN40zc8ExG9GKowtezNqp
w5nP4fUABewrFoIk6rXTBFxzHWySlkCMkTPE4KAfwaDlLxE5IV56EO8gdEZ0NrHRVO+2nLU6E+OF
Xw4hLb7O2oW/LZFuWXKuVYeLZFOeisccjt4mYyR3tls83YG1v4ZF2CVjIKA311hl6xAErHBSSnqq
RO7VOVDPe9gujlRG0oyUzalCxoWySWhFOmARYyG887Q88cXfn7RG8yxUSnZvLA2OhSsc18pSytil
6oiwDJfEoSYM44thGPSJVC/GEjYulYyMAYiOoPw+Cp5kaKQTaSxWA77fsiaxsQooCBACOOJv3Ptj
EJQjXunsPQtjEGiKaNFV2hE89FpeZJQxEAuVgvsgPVx+ZuWgUP5FHOHvg0zvntZgyn1aPHhvpguu
VBpCOZoDXXiAMw69B+/NwL4oqOth2iw0zFGYVAEFpD3D8cgwW6IFf9xNVQynW4TdRlZwl4eELiju
WjeWlpZKqCnWYjZuOrtR3e0Ln9zcUaGZuryV30gE7ByZgbBLNPz7IlfPMyN+8vcOk0j8JbuU6gPQ
WEhMXQtIBpjyUzAlYl94lC/lgQYzWNf90xtc9O8fK1IK2ns5ANAfRlOwhQDjCIsCFsuVOD6dsG0u
B30/TJBG7m0l35NDm/2ltzsYtOQgaabngu1KJbWAsDhvA041pQxUs+PddLBN5cAOGsXqk6P3QwT2
lWicdz8ZuJZVlQgN+S2xIYkpSULj2pfdKolXjFOf/TLgfFTVUgRvs2EgaTLyN+3SQdTqk50hbqFp
FUfVUyF27tOZlDx0P7jnPUImyes6YpG7u0VjGR8SlGReo4C8PAxcSxreTxUFi7rbUXSHdAwHXslA
gatr+XKLh8ZqIvv7X5zAl8oIFUtOAJ+1o1t71dBVBVeFplEKclbjpo7cFnmBKSlRkMwKLj9bhkTC
bRflWS9l3gTmnrPjBi0LZW0umyNZkd5ymDJNhX1FtnMyA0wYuI0gtmPwCnRlV+88pdCKj4DD557w
ogetL1HRwlL/pUa2LKwwrbsT+WN2YIsLEnS/fn2oIzuoAQ6mGRdrcSLAlTd0xHB0VEXhbxiD+u93
Sr3LlawrhNA6sxhrzQVaVJPW1+tYU1DKuDOXh3vDPnsno3BrwGc/zwjuaeS1ZX9AVbyRL5Gcprqq
sKQSZ/FrSb7tCym+zx8OaHGNWVcvJaWPZ4+2OLSbna9bur4uWnCXV40319vZJmxroV8GkilBtxP7
Dd5KtYTG1mhVJxMJMAYnu6EI56QvlJMS1qEfA8EiQwK70I2PnVP/F8gNUy5+A/lH7zH8JtsPYUNB
9FBRN3A0hpcu/6DrQ7E3D2IHvZey9ETO/A4FE19wl2yScoiPxLk0aCzVeU8bbnpsDD793Hw4kGFT
BFvdUVVN7fFMfuGG5HNdcg6WgWBYZ0dZFgyRkpc11BMKaQWnr3HCYr9cXORn5f3+eSjJG/LQxem0
Zv0rTVp+IPfVSEpJn1VMIxiJrpyXlLHbcV+Vv4Iw/yQxf9zOaiWBcH5M0D1FDgs3/NVLqHl1s2yR
KE+WsLELilGqZYiZSTdWXnUGTKHFFTwKQNZFlGYaGahRW9oQ5nFw4LgSXkSUY98/4Stl4SILF6ER
tCadb+DLFzF+vkr6/9YC7Jela1S3YS3An5+zqydSTcojravLROOPRTj2m6rZDGySD/XpKxBru+Yb
DY0iCCeFr+qZewxl3viN9VpyY3+cOGVedwnwZ4bjAMV0/2RI59147OwNOXN+bQmOINgFt/6Fs26J
8LqJRG0q98wMakj7twm8I6lAEENJdST4/Tb/5MRqrCpqBERhnB0ls2zUDxBJoWh5j4T//CwTFeyG
PqmFYIdd5erMZHumoZ8yZ1umfwlaaR1D7GPasz/+umvLwJl8qSIPsfzeXspvE4slgOlSe89xzYaX
4eGE8OZtXJ985Dks9YKx3S5y/5Ep83sR3QLwUyEGVC2JRzMP12dsn7baLrI0hKCk+IJjGSmx0lUr
oigkAuR1q69DN7T6w9KIciZPB5Yxzo7FucFKwc77bkQM2BPqh9XttqOuRh/pf3vMDNcrAS1RjYs4
uBtlf9pYpLd5UxxgYHJWozrxaeEwd55iw6JQnabcoYjgFAGWp1e9cZaE3B2t3odgrmJv3wpqCON+
H795MPpqevSQCbKdXHzyiJe+1xk01d9w2zArsbDaieLTBeBNsIXrpw4xsUnDxPIDgAs0TnMKpbQf
Eva9Jn1md7bc8uzHuDHZDp9WnmhQ92aQQ/02yQkqA1N3w0UbjpanOqgASzoukpmucIX4YMtMGy5v
gbQPohJ2OWCWGkwdl1G5GGGlXmVVHC2LFCNOEWll1IETWEicaq7X84bW65k8kQ52AQdKRYj8Tqw1
n8j4jRj2MTxEsZGHwChEnDsSq7hcgKWXLaaYcG+nJUfrZsck6LrlY76vgaSFYHxOuWTbtFilirgW
rwmYTcx57/VTteoybqC63W4QiiTQnT6z9Re/CqPN33NL7+T0ggsUVTxgumKYFvW1cLL+M3ANmTOg
6H3XSLjnOlaMhZpbzzyVOPMYkf8euBXnyqz54AZ5MKdefBMtJP+Sv7dHAADVAiBdr9hJx7g8euAi
VaxSUjZFkM1wKivWgt5Mvm22q5Ypx+TkJefIbGqEEw7zjjzuHIluU6gj/ZpzdE2mkuNO4te3aJw1
9IkNnJHyGLSCRKBtFFURgN/KKb0RVnilA1BPLUaXMCeKfreqTLr7k//JQPuXw4WmkfhUS3LSPBy0
3oICGDHFSifzmgBEqnffzDi8qb/A6pPl20ovS1VJQuHg5g42/zOucZAN1s5+aJPb1FnxgTHS+ttH
cLeU9B6z5d0WCn6au5RsNmtI6zPnqAmesghu1s7ryDLzpnaPVtlOpbK9rTbizy0ggc2IPsuAmH+K
h4gc7gYVHHgLSG2jDia3VzckjExrxFnLlPYlZmXFWe5DA3eAnB0K+xxxspg7+z2zNaveDf16sZ6I
F+KJBG2sG8Pu2ArObUYsSMdSszgA2AoKPNPqjspfGiTV5FXcB4asBZLYJ/wqDMQDZ8FgmpHUPyCD
An7PEUUgFgo4rOCZ/stZSCjDS24dxm3+H6lNxTn9RMv11qbIWHuGdV5bEAOq9d3crKkS7DwLWzKb
nr7Ua6LL8wZa+ejPmi75vb6fIIAtIfTHQ0xMA2m8xxbikuLpFpoEFOUyrBtCsMD+YOuisxVMKQuN
Q2/LiCQSAv3zpVdANZM+4cL2kfGx4vh4PA01wz26H8hGdyVQq0NY5D9F+ZFE7R88RtkKrriOPrQw
ZMiF8KvIGOsylbPO48LFyx0N+RxfuPgz2qMAr6DnSX8dfwEz9Z9tOpF3e4Rb2tDziC64mwew0rha
Y8sT2WT6k4AoAnSWxfj+th/j9EI4SdBMsNTxa3fFKoVtrHq8wf8shL+qb/gfGv9GBKo+JeK2vRP+
kStiJxHzsGLFFt10EjTTpvDndV1Mmt+XpD+X4vV887SOEiIVoOsOISG/tFNvsQLxmPaZEUXfOcm1
z0eYnIORJaJ9YQ21AjhdYXp48krqRyRPGpvAA5498WYCiPh8bxLQ0LHJ/spuSr7/EJPGVfpY00l9
YChw3IvgZDDO6gGqXYadTvDRNKibbCnDBzm+SEzoVq8QSCdUv5VqMQ2ta66HoIT2Wus++9vSpcMl
Uj/+YuMedHXBo8tD4fbJBaPchOfbmtG4eFvT+vveZ7bXCy4RoPVfYd+nHl6I/Ov+rEx/BJ5afpW9
Ud+Bhl6BwRmIzu0OtE618fAjxBZS0v5GJdOcM8o7kmIAVUmivMHeEG3/oAdvS8DW5BwSDkWFRwSJ
qrKlyffPS78zOUn0qtLc8JPb3qRt9QHNAcHBjR0gqo0mD03rU31t/I6R+6yLfGaxNuVwU4SylDeP
uuj74V3XiUPU4xK+ioj+UfNWwsSuV1aSte40h7T4AngRJwCAOX3ZJDpASbCawrBj0vS4aT54pkE+
Bta6dXUdxqIZsYWExTN0w+EgQ74cwc/YTbqClO6uqXlp4+HKK8cSpbYyZ2RNtVbA2cFZeJmEGGtC
KGWuAQKz+pBcaXSiDhDtkiDADAzUhnbG4uYRsP6d23URH4XmobBG4KQhLj63lVkP14bDlYfxz7Ox
6VMRyLQEn3hXckkjvFnl1oJ9phM3U62P22KNkFkWrKVxf/QgfoiaPAP5kqvfwyu/nhgtE2pGep2x
xMRGsQE665qvnyHH4WPJ+cZJ5uWvASI0VbVm9eKNPb++VB31IhtkJ4KMQMLJWjjscVa3j9mMMN/B
bdN1kZO5fIcPKqPktq7uDHofZz5JkJOOSoj04E9vUJEi+ctx6tJ/VhfrYaK3QPey4IoOYBDlYe/m
7mlbhdqUDOm5qTSKGmBi523+XIsaysiHNz7vv4idL5r4cQzuSrYnaXVTh0YBqwbggptKIl4q7xO5
KHPClwPfQO/uJOUoyUKBzui/AB3de+PiBbZE8byWGELR0kXfBwhriE5mvQa68WB6PNcoFAF0wkB9
FJEebG86/NVYnILfsOuIJXvNXybRCRIft+xhJ0MEaz8PS8FiR4lt6pI6ieWW3cdh2XVWzBx/71eh
TA72vlM2+LBepPI6vY4twAOw/d2IYoLuWmFoYHOzVBu7jL9z8Si8haqOm+PCPqylCW3ckxE8eTLz
QnGzDteukOi8SMisIog6+j6uSu+LkSRTY7FSxytf0a456qM+K8kvmlizyiTDLZ58IAlM/1tEhQ/i
ef0DFhWLly4zX9Sv7sphlMMFBeVeFRSog7emRgAI6mln/3aA1ACWgrKG2mT/BWGBhA9uLBBpYgMC
CFGRbtDDbKxONCdRNPwTN8eoR7AlYuuGCLx5mxGfjcih0hS59WOAeNesDrKfIIcfg+hbtD01PejR
hI518Guo9bHHa3GlhDPy2riRd2lSsvEgEMPz6Qgkglwc2VC3pTqt1eJotGFg7YahrF/sGmGyOrnS
RP4x3iYFGE5pl9aHmtAGt4yZSNDZ4NcaBAlkvafUhs2fZfPqMWgrtRqzMVkpiX1RTRePhgCwwJOQ
siRJ9kwVrAk7XSE/WZkQ9/5BRwGQKrqiqAnqwbMP8KQuOW8ieFI6wDixVttYxwZ/8vW1oHhhqC6x
5v41/9dIzY4sMuSRXutKSkW0IFNry4Ew7tD22olUqLBtBQ+wTuBn+HMeJieb3fhUlEuUS2BY+S+a
z3AR2XVYAJAislkkrK3VouuodzU/yTDL3tooj2it/no1jmuQwBDprqHrMlUCBi02xHwSU8YEgw6y
AfRbI6xzz9JaqyaU/vwfXg5c3QM43LuesbAIjrY577Ji3qlyvUtM7PFaDE0iNOCSnt1iweCFUj2+
98Y7f5bMw/hyjqbBvMoBpGKR0ChPzrZ6kt6zByqI+jIulVBOOhmbSeC5HxPh2i070wiQx6rvOXof
dugy0ekOAjMNZ+hRkuKoBmwhzP7WTGnMOXnFZnM3lW3DnK/gYIY+3/fWAroEtnhw5qK/q4aEYbsP
uqBxHUGkIw5zI4UnYr+rCr6SbupyDYwRg8JHomhUwKxz92J8hETDmZbwLEccrWH6pambc1mHGhC9
DRAali0WpBUUKhLYQ2y3w7rPR2MG5SS7M+Zb9bVt+VcOpp4kjQM2sRbHIZDd5XcVuGE99I9UZfR6
wV8QjMCzzfUsRrnCtnC71TZGapN07AFNFJXa1iWz97IDvNg1nA5P7ExeOkBoS78cVZsXMhyzpuAn
fNMdKZEYOrioPN5zunTYTFrClUKGrITz9R5QlyLvr8rMt2AqaB5aEYUh1fMb5yK/EKVYMTjhTrFI
it/8A4aqBrwIMOlFGifAOvXWY91uojFd4Fvw7eMo4VSq0FdmaLLDXBN6nV+LFAuXdhhuxuMoj+Vm
TKOiEtk3LQsT+bKu1+GUd2wT/mvOg1ee95Ao1hqqiF4XASw5pom0I7WbrVGbspLch03xOn/6ylXz
Lu7Mlc9iHaI1M6wyb5JipBZ/ygOo5UNEoGnVSX8dWs0KH9P0cRCLiXnAN9X2zpUaVvPyoL0MXggH
WggkG3hxO970YpncSNfQPkLsfipy5ADDmC/BtgvJT9tri99VjTYWRcC6MJ8fV/rqwzBTCV9x8ZyQ
gDIRkUxpUQVdJbNwmWzU+Sc753PGxjMu99tU7h9YfXXhBPrQr10/Byb1N5vJzmuA/KKK5XZMO4by
vvdKfr46SE03POfjSsIB1NpaYPkPuMHGs5CfH/4jDnOvZ4ML5dc4WEwun7PrWgpEJSnwEcwT2pk+
VDgM4TtV4XkVjrfuwjaGP/NIwA3LmF5P0WghHVNfVXbi4ZE+SD4ROa0a6rsocuqiTqvUyZxLfLXt
iEymvKmyj/XXiCXydd8DB/aiAwm1uP0aviltABf3qohpRMRavb/IWoFmEf9JsRktf/pWDtzGqUqd
L++/CQ4yfvDSCc4m2s+brEOIY6wNoD9kT0f8JLzYLRHBh4ws+m/w7fiOWIH+wNPjQk7Vg+F44DX6
pm8f24/UUnZIUJz8uOY/S+lzhp+7w5STvcZoo9U2dyyGVa9VnRZsIBQXhzk2ci6j7/ZgJm8HtBFK
S8X7GiZB7rTNo85x4VVnbuun5kjcxbkCQT4HxcCipVMYt50M0EVyGdu+C1w5NHv4bae4WibZYt2D
o0BP8KmyL2Sv73Fo9I3gMvf9DP4Q2PhSYvHcEMKnqIyWm27COB10VXGrHM1BZTjIpv320gcm5z35
Pn1bSA5ZUwKfB/pCS3jlsghp6/CS8Ru4/+jsyWnSpm1ayJD4t0rp2Z0OPt03aUTGmTeB/hlSIiNX
Gw7ehjkW31HZ2RVDlJnoskteEz/5BPvrJOowEkmeuAs1yudteTXYShP+M77G8QeOQ2ZQDSRxLTaG
Lbe4pmci6nEAUj7wx21mLR696DN2+Ih2kCFmDbhlDxaCWEg9AVMq/c9mFiQNo4z4pJ8DA9qcvnEt
PxkzG/ydg0JixrzoMBSs7d+loKt2v8Z8kWVu7Dyw5l6dwH743cjHqOkiUhtqJ/+T+hxu5r4lje8r
W44p+P0hdXKQlw1e7enax8gLJQKXYkWlM7HnZyf3E58OBH7HENpdE30Lo6Mtf/D2vW5OZOs41q6g
2XIobUt5yPkGuXTOrpiwMJO7BjdrMitlTI9uhnsxpt5TthWcqoHiICgIKRdime+OzKFdRVgTzeYO
zUCfCuCn/dT7KgKWU65ZgPGOQcRqDp9TQmmWDx7yKpShkmifZEtJOx+gUd0AbgXUXsCzbWUPjMt0
jIP5u/GFpkM2igEKmPmIqqY+5VMrTXMwp452KwdlEZ0qvVGNa97kmyGcGYjG3kZYRFlsdQUPa5T/
cNfUVbgtIjf6LttQHSKDYPAubyB/zKVpFVlYCJwo4KA0Y9Bx/NkrVftpj7JdidJSB+tZNo2xR25V
aYtIoUh7wEvbzkH8nv3uEuT6KMy6Qq5koDDbyD2puc6vSIv8z8xNPrI2CHy28c+2tfaMKlUXPtLL
bbpXs+5VETjPl0eV8nGNp1KFVGDEGZclewo/EJK1eIZZ9/2bMoZHpH0rdlD/0zC1I9EfN6nPJz/x
+lcPNx6c5gt1seea1OrhQzISkT9qjaJ1cjEzrXgE2vI5Ch49ZrR2yCpGQSHgeStIu6OlIY1/wu8u
rCD781wKt+Ik1H5r4qOatCiMt/+Clu2JqlHZ+vVW2NMKaaM6Fg0MRJsYqfVWFMe/8QxyEuESq0zR
ePEHAzJ22XFIPgVEoYYArM1aJwuUZQaxpaonBT92sLyub8p95OZCWuFtbs/6exo5GGyH8neOcqOC
eWr2X+2CCHE6E45wISmhKe0C1qETxTqvUwGwk5TpsW7wsyksdlSOnlxTSqige4nRWKgtt28nkRWP
B7BiLuyK+LFTAVjFZar0mkoPXBfmHVgnpCaR7ZUKwPGOuvTBveQGes0IuEaqVtGvEoWlkEFAREuf
c6K4P5Ut99qxj62VckCjeVZCg9aXPYIvWpAMyMPaLGRVtKLsr6teuPVg1toVfImQ+LOqnUQD6KJr
CBQ7NOEf+mXiSUj8uvOiPsN69aNTZnxZzm7JB+XgasnnsgJZVYzPJReaOgxinvy8/ZdTiIxz7YUi
oTfP/cLNH5IqHxTkLIGVSDyixpfg/9/GMnoAfysbxJnIOYdwrAWa5isqNUHmJVWs/fcNDsrag2fx
dSJUdIOh0DLmhuSw4I5qpmAzS9l8SmOp82YHrVwpyw/0BwLVwl3uLPb+8mBx9ZwOcLAHsbC73uDD
xa8PkPaeVz5A+l6OHHIHa6xHuApICmhK7785sdz4rNpYM7hUPU8G89qB6fhy5Wg7LKFcXDJsd4JM
/M3tYmtFR7Wr/4He69YjSeygPe0JmkbWY5EWvQp4c7JOHH/Wf7jp14uEAKqN1NHaX2M0pXmGPaVx
nCOwoDeBTUB633vP6KtwOqhKBASRg+aFcr98yz50HJTa2XhgunfRLMEbuzUZzD2qoN2mv5nbbFkv
Fv3jKKQP3FiLCka7EYHgHbz/0kDT7RIzhrJCs4l+ioEHj6B+twuMzr1WFaGBasLaG5QAnvKgOLzp
el5GNULNZxzkqYtsbv+L61WTlwaSjIiAc/IGuehzLcWIMbMM6242RSsUuG02zMxJijLCD7SCSV1g
/wHKGFEJ+F9NRavSFru87dYs6ujBzTIk5UuDVefFdVhGacj9mG0d10TSh1WRWtY+B04zRbju8riW
eG2Yfwm1uV4/+5MD6wwJUIbwMvMlYwYvib22gZz6oTQAK1w6PThV1NLeV4xiZ4SEH5ig7xYSY8Ni
lIfx3X6XbpciznX+kcGVRMk/wDa9AkVfd8qMV6sIqQpvuCrCeFOs97rGSD3++UgnsCxTh/L8qYwq
NB0SJxU30le0LnPlwUq6xoGkeS3nN57e/w1fjZWzGhmfkIOAfD8/8imsDce8Z7Z5D0VpPameVIam
pbN2WE3P23voOPHeafJJ5o2iF6/QGDtfBi/8P3r7EJnkrPExB+uIWR8aNHh/+RQNUnla3oUlbcdY
2lg6+k3280Cc6AwioUTgyq4zT/EhnxStJ8JnL71RNAtYb5iPjRft/I2j52hl0QqMnc6IYroddJGE
XzY5jZyUyG9sOakoj1QPdzBcOLDyVQQDYKEYPdMfPA75+2jnr7qlTkvoG5pWQSR0oGqGYWdaTDJ+
v8x6hrrlCZE39Im39vDjwrdQq7XhYDv1GzzjC+/TCVPHSszjerXln0GFHTQ4jhLtC3SaAKJ002N0
WVkT66wC0B+NlPOZgK8HGsVSg9lzNbIL4iaFlWMIt1wD+vfoSE4Xe+W+5LT+4lBGNvhDgmnQcHh2
F1WsxU28Nrk10FdqBV+uLNrlVDMNFtTOXxI4hnFSVAuccBgYhPz5/aNbIYeeTq4rOA+D3LRPxCuZ
MuySGbU+d7wQ8Z+Fx8WHYwC9DwMMDBWPfJAdvssvfZQqkablMP/g1nJoPdPAsv30CfCH5em17mnP
X6VlGN9vwu9o3BalFw0WWDP9yGmIh+UowraodrWgLe+DRe0hQQoI8gmBztC8i6uq4OcpLPAFW79f
gaP8TJCcAjyC1vQHKKirQB0/zZuGdT1joTpakfUZTkg1j59ZW0R45eqcmtteN0jyFM14ju2TD81S
cQapETwD1R3r55CeTtixHVMVK99uNWJdRbVRbKFReZYOLpG0hlWITcEJGJA3B35GXjd5uBIWBQ72
pc3YsVxYmaZskbaerkkCGn2Epuachmg+oPw09KD3+W8d1GNmgItVMvI+OX//sA9TG76Z3s57rYxi
T5qw/C+B/505bokktH9rQcoyY4YJjemVWNYzcq3j88UGZvp/0avmp7RvF60XxgTEhdMMEFzV0YOy
GqQUveA6FbB0DTMoEqRC2wrASn+sh3vr7nTsNYwyWPxdnuNfIzxcwLtNK42xs+ALTxjlw5jx2sBw
oDkxRcvJCp5PDQbI7md2UVTgDY7rFDxpwGNmemHSN5n2cfZBQikztdzlHi7qKM9ZkLTZO7EB9u5n
OgcfWm08rQ679xucRiLieskQBJIqFD4jECSrpJvWbhuojOX3S497bf1ZBUza3zHffKlBW9FtM5v7
NW8PCtGKKLI5TT2bONyQH9+5YLT9lXvlDXnGuu26jjzo+rekGeqq2rriSRtpHuAjvSYKgMbS1DNn
uHJ8XLD3QvBpoQlKfTPrscmlP7AEnjsPLnE4JUsHEpcgFSJOjjIO34YhBZj8Pgn/qMOYkt1FJaOw
QnUz6rTHrII0Xv/PKE8yxL7K14EvMqiEBrbKGS+IKD6QKzTAjX9QFcttcf3NkpVr5uoUi5UMTIu+
TLW17tVGoeX7jXn5KbIwDQddwcZPIpoTv/qd+N+fKOt/Ac6basVCjgGifPjYv+SUtnxRAemHq47E
h99MXbd44a0JQJn4nWEsnpqo6yFs5NgYIwPH2Lf5QrQtEDk2jcz+hsOoAabFiPyXfJkrEljM/klC
3jUPg+Hinhe349jfuLr2GsCZ4NsRbnBC7Oh8qUySYAShl0wntyHdH8wk8R2XspuSS8JSlNFnBrug
U4aAgCyjc6I4AP4AnX2PejcXEc1uX0fm64okTSZhK8pRHXT3Mn0rUGS8XORUAM38SHLKU2UGkn0d
uqba9vTBzFpQshs4ApxO++IUiPUJlEJDbFal9oI0zY59bpiPyou7D7iIdAS4v+6RnsTmK5naw+u9
95y4yRkCd0Lir98RBs6hrANnfT/+tJN4TVuaSpxKlQGc0IEkhsYpQwnL8yiPbnWcB+MEzNAb8iwv
IqqsOhtPiiYkezco/0qKPei7t3iXyIFGJqlHv9Gh1ijWKxHw6qEDKNJKfl6OLPZkZemWUqFpofYT
L+47YatO55pxXJtMmpxCuhyMB1c0xS0yuHGO3pgYP1uDGQqS9SdxcFoCwdfMZfJqcAPs3y1GgLnI
Sj6tLKt8BXqOxc+NIsqldO6CYb5eTZQ9xWX/WyafgNBIQ4oaC+tXBAgCTk+31g/CmoipjYe44qhd
OhW0XykL36s5B9q7pg/WXGoVSCUhgLnlyeOhskSy0D9DHyuXQlOvDef2uYkwsYpVslrolyp+aaFn
QevYa/AE+X6JBZiaB2yKmsWdUR7A22ZRaD0tMuN461xaT2RX0m6lLRYNRpfBH4IHKvzHmSlt7Way
4M4hNWSesNzNfEoGX2PVCeUu03AFlt83aigAr9Ezu/wSUEsrY+LTUEKxcJSelrfPSvsx0W4q1GAe
CZDz7YYw0A78zRWYT7liy1JLvAGgr8A/WwCN1eAYMvdiZtyHxyn93N7NfbaJR3YezESvuPEzWRSF
zYzCxTq42o99YNxGehPkINgCqN1wtzEqAVBpmVuqELT6SHYn8rRgzC9fFy9DzuPOTphgVDDFWUyZ
cGtbKQH8JAC9u1GbQ0CQTc7EadQyIF0Q69PrOCcVl73DPWHIkpJ1sjH7U9yutxZDLuk8qbFYEZU1
LCpWVctDW9QtP09rOkugJcWlPV1i0ueMRqoJTeKfokmFtUTpX7V8Jq/eduYZQhob6w7MypjrYCcl
11k5D+INZUzQvE7B4/yxlKZdnWg97+kzPMBt7uCj9rcbiOB2Fp+ql337/p46jWx5fpiugNhPEWX/
GxOFLVpSDZI2a6dk3seg+R4sjTc1NifOtEqPDnRs/tFtzni5CII/GQAzXGNNRbH+0C5KHKVDNleo
kO6Dl3d+6xWB6JamrGvxiryp+94stVawvuqRv0Feuxddh+dkAyN6arS9MUxB2ui6U+p2xISaz67S
0Ivio6isqPuImO/I1k+7EXVRF1G1aq1k71a+C/ZKXiAN/cX2LOFk3hYBVkejmnWDADu/8VWvrgmv
PYMM3uufrwxDvmebC+sGngTFy+b6g2c2UdHlh+t7CMsleUMMno5aATMWmukuLN4HyvSlrc7ow9TM
0pBylYCDp9TybteXn4euhKoV3qA9XAwyQy8DRL/6OC5hq1Lil83acKCf5/qBeE9wUdVRoai7R85T
H7uhnk0MuNRwPUdwU4LVo3M7IwZKUp1xrc7WsY4Wo5DhOoGysG1P3VBH08hMAnVI38gadO5aewSa
vqU51wS35ClJwM/abwvRLt9jpio+lsX1aUNwN3LP7peg1ji3kasvOEegNtNBu3HmAjZg+qZv+kGN
6KQh8RY+ATSGTxAPVpqMFQdE3s78ppLrOZV46e9l1leVoDApGNYdYUwJlKDXuR2m16DMNXJz3Yod
c8ifWAOpuxeiXF+Je84uYUA2OUeC6kC4V8bKxUJzZgy3Zwyi83/0MNnTXTu1jENixOkH17sX0i6C
fXtAFEB8Gph6WA9wkIn0Iw6Ctks9kVtjVHpSDF62Au2jTnB7ukifnP3wpMgCYBRxQkrgDI3uSwt5
hkPerbDhjT3X9BmquYiSlt98ahYQQotl5uqf8eFWKMo3HvFwDALfWy70VFykH6rCM2LHz2+bZNy9
ZHTBwY0aec51PIjkPz1ITdiIhoersJJ3iNoQa0WaHOA6XubGWW1q8zPr6adp4U0KkHDOn+GQ6NL4
CBL/kaWeVI6oVhsX4LWjVhX9qRgA81sIObS5fIdaxfS7BIh1DqKMBWcVM8hcztD7VYX6vKQ8wOgA
BLwZCFxSe6my7GXBgqKJb0XKzRBbXeHrfQMspQqlm51GVcT7T6o7mjvOya1njIB8jJdD3TipmJn7
a1zAKvYt34kne3lO9m9Hhl0Q1mbQfgsWfjhvbHv5NYJHF9XaIxE8FVKWvOAXObV1EDDFpUit+ANK
Uc1TQj8JNmp9io4Tr2AwVG2XohHICxayVWBWJFtM1tIYDsnnNEn0qc64dlM1UM+j5h/pWGMBbaaK
N9OfS085gqxN7V9K4w/RSCyKvv89i9VVgCp1+yePyIa2X/IKuyNA2R7dKX34Hf1RvS1JDOpY82GI
M72/xsdYqf/zB5NvWYTpS/KjyGnJMTYobsDBx2JJN0nIuNBHU1jw/fLQsrni4yqooQ54qWcbm59V
y33AlL2RhpA22UR1L4VevCOKQkcbI1mf3tuTXZ50LaTaUFrSg7IzNXcCt55M0qGLBkJ6/FJvrkYj
1EZRFb7iBHrev3DekLFT1FaXAruwLO+YMPVMRq0uPZFO3aPUEbdV8zDBSqVmBxMO1RA9NoBqN5XL
kgxlyiKR4xQnQKMBz+ie9+ZgNhE2U0KLCOCZ7OJEF7y+PXbcPAY6kgDL/TtWfqzsJcMTHj/Bb8KU
ku2V4VoqmWqeJJ3GWfQhYKco02jDMQTVRljARH5UoIxAy07LesWhy7l3JZ+m/80sZEIoKMHD0FQG
eEcA5TxfiibURGwE0oy7uN70IBTfAT9m9/HxpvkXAhY0S1iorNzXmTg4fV5fdCnQiLFmlOdtEcMY
iluKVKYHXcucF7HeI1hhU/w7xkQPyVuO4EFT9cjHwa3ydCgjZqY2YXlSmp3oGQtIKESSyJQENIKn
YadIBQsExYvdGVk/csTWPZNKbPmINsR2r2tIUlhXi+Sg0mroVfoAH4JtsxO9piTZNPLmwwfs+by4
bdxgR+xLUn3KZCFKH5iZhbZtOLUhFjSd9QfGtapd6mWpQQz9SQQiLXb02XmOPgyXY1teST2KnxfA
rd0ACGg+wsYWJuDrrnFExS69zdkIbcVxReSug3rlEB+BWNHV2cOJANabjTyQ6KFT07qWnVhLvAwo
Jil3oieAL9B7N5B3I9E15hagTL9Zp/F1Rg8oLllrNZGNZjssp2PAMLhcstlHAJWbMzJYNufmK3Ya
i7qaKJ+HobS8QGZVx0mMBixGn5a9EgzcqYwbZLW4GhqvGWs+stUW89FAGkEobH3KHUKiQwyRRfKj
i3xDqqfmUFA8jeZygDGIlgmB7+z2l98r3j0J1S7ygZMMAznnPty0x+a9E7t8lJUx2LGjuSAUOvfw
x/DGkrcaS2OzFDYm3Ny/MjI8RjFutSVxIPHwPThIK3zKVJnzwlzmP0jxSGJb0nltB06ZdUJqUvZ0
R7Ppz1j5gHYswksNQ4OBwbR3CKiA/yhFhxtbQAjtO/Ix/mdxEDfiAGa1DrJEFOH1MKwRQp47ipNm
cPRmKWvcqazBJptkegwkJvRMH/H65CTDfQpzM9+zyecUI0uKAH6+stizRQ7fmMzAeHm/Oys16WLp
K9h2bXnz0GrV2cX5EAy2NeYyXoJJJFwkquqIF8whU1YeLVKcqN6vUsSXNYSba8ImU5ewTl534gl3
8mkfhJcnkzbmSo7gnOiq+gytNP0Og1T2CLGCFODzGwYHObAJR1CfX4JNhnarjdafzUejSTjnuf5u
s3Uz7A8yXKApk3LPo9ZrXT/7OJyknmzEChnZbZQ1QMNd860OoNUH6NdbkMkMazZXuH1Mk0TBIIYh
9eNAvBp5ezrUvfkyPICnXY4GgAgJn0TFkBM/Z4c6R9ovyPe7Wuf24cW+ScVghnrCXbyzMBU0NqYC
RTPTeyCkiPU1rJKVJEwfMEjHtBjr11dgjvo1fefVB9jGesRpQ1TMOv0HdD8aK9CWm7l7ZCOgSTwl
CidsqDVHnGjBcDJi40Ka9IF8+KjG4XXgwQG+kAxk78g9b1d6GvmCJVXzhEgSoHliLKJ4Z89DkKx0
3Ejo7cO3S6aUZbCFTMy5axVnZtMUsPCHrFwHZVwTlYdwzQnTgxXHEHs5hQhdD/7c9usBBry4VH7i
eHrW6+pn9tzFdVFF98MHjt9tfjrjjN/sW98IdQz9vxLCuN708JbqglnQ/zfXl/yKftOemmDcduwm
th+px/8riIuPczEPRjelK9reshfJv5IALomRMvf0Y25ql2zK4GcHB08bSEB282EHE7bUi4jUu6MA
QFclbZa1S5HHF3mbdmCSP7pKlGPAR/hEqvtgS1hPcMjSUkfz47Sv2o3jvT5M5MEIe7kttpQmWZby
xgoxxkMIPElKkpcyRk0y4oNFf25C/RvgU13u/aKyi63GZ5ghsAy90GDGGCY4PrDl72Yij/dB5K36
5Gi5SSHW3Pvxw8VbzOfhi8htcKLwk7HiKVgpS9XV/aLxxT8kut4TT1Yl36cXYtkKv/8VkN+IshTe
ZcA3dZ47QuAFTkZgYe0mkdKmnfobVAfIu3Vg+pdEc09O8VrfDOfPsgME3ycXGVz3fJTyyszhTnY6
dF7lZ5GggXsPF3+WGwEgmu1KHeIo3NfYTDGPHgXWWL56dYQfN3p7z4+4Fg9T+gmSE2mbewwTX69i
OQWbYXQna7Mcq+qbBvIFAQLupZnRp063QduKmgeDkgCHCcnEIKiZ1gYNdqyX7XsBXH/irrVUV3mb
75phUYf7PSgl+SCXqp7wFlon+noYicWPLIVmJAjx0FooTB+zNenzCti8cpRCDpz4ZlAL6gfvHXsD
8caHb+cuZ1e61Nb7rLNwL4wR1MqgfgENpW9ex6ghPvwf211tXi5cUT+Btb7dmj9v3ALQo5Ey70u1
TBKinuFvR64Gsx8iDwS5J+Wy8isjvKTB7e7jalAQKsBxC9K2zx/aoyoBDCiYuFWCMxDxc9JhTuKm
+vcObdGHmwHPj+YkHfw7Cqrov7Z2DB1x944gHu0sHVDS9gApd89i7yyxSQR4KwzSn2Vd52kw2JYU
T53JS8TGx3tZQoNsriCslndFZc8RxcZIIKTG2p+lCMRocaQX9mAULRxn8bL4skj8efvas+9tE/Dr
6NmBsG9EPy4XIeX8e+iQsjhlgLyTZiJ2dldTNIr59AoxAl+dFNYqdY+VeVlDQN+RYm+C6+gfW2z2
993xdlLyw4fCxtBleGPwjSFzD5qGGQwAxoorbQYLoeEGiwJ3wtiAvNkvT0Or3sEsbca86C0H2YSA
n3QrOV8RNdKhfPwyAhHM4uq1AtK9Ena3TmlAOj2XusMEvDnvIs/kxVg9zZLLHZtWqZNLxlqroqP9
YyaRe0VbIrNMKUqLjHvxbg+s7JraFFuyYjnYpjGJI27bdTQ4lestSdQ7adYnnnSmwC1zp/VRc8r/
cnslu2ikX5KKynAtYhNUcoU+GMqVbnfDRQMmjlRhoe6zmGW1wqroUrlZGUl5CEDyMfcyMjbVmljA
OkXxrjLqaWxEb4T4vuiAkmMqx1z4jzCS55V5lUTuL4ABObp3DdPnilVhTzlHgpHuOSM5aoShsj0+
4I65y4LFAg83hA47k2ekbcUdWtMnSMZGTBACpdteOtu7L0h/UUnlt3asZoXD4APZaddFZAxiaZVY
Ckefd28Im/9i4ioKjRFFoWj8kV16fMP9GNQqADfSaXVbDzH+GsHzlzY6Z5IkiEgW2lArn9JXxxni
TslHWgj0yZvzuY0hK5N1r1IYcNhV/QU2VR8hhgOTbpUWvhp8USzTeWir3wp9Dp3lnwtO2pmvrdib
+OgvBWE+bi/T6IW5mVyy/UX2qs5JjipyoTQDUBbfruNy8JUCxj52xr2gqWPO5R8FmCU0zaVO0mes
y+3SMsFUoKjasScEX7ggWHlnpqV3cs5s6fiFHgLNfO2YmPI0bBHqJmiuFu+3iMLAqK2SvA/46edH
7p9pAxNA45rMaTPcPBzRR+j9FcVRsWB+5NXnP7lEfQQbTwF7fGUD+B7hZFlZWjNml03MQgKVh/6/
OxQk12qW2HryT3lsDU4E8bygrN9NOpAjDodfzdICVthGyy6qoH2FJYcInOoAfe9zGOaezXoXDpkH
ss9tMG+MzL4Im4SwSGbiFKDyDg8iNNqR6ii82FeCMUX0mrGQSMxiFiDPUgnU1J+jqEli5DSaT28Z
UuerTq6r7txapR6bhSLvQQIU4C8di9AfgU0LnaotFqXtWSKSQ4RFN3a8h0W6qnALYviZoUZaTHbk
F8NNYjDuzYwyyXLoBiv5dD/qI9GAu5HiynPoSTIi8AHilWxfJ45/1MLskmF84jHXcRgoEeGWwLIs
WDvnCyJdeKNG8U390tYv0SIxgFpPmV4WTNNMQFcyuptziO332dSQSWOuVeC0jtDYhYzWzVkuRnf8
uXJ9rYQ31HVZWT8q3raJ6SftHGKeVB6LF+45Nrj9tnBrlGDspOx+yyrZbF19qq6Dnn5+TuH1m397
mcOKc8e5FtGvMCw/4gfukoq07dhJiZ0mj4mmN0cczFRP6u84ZpslzjQZOgcstAmcrWYPnS9jauYa
xB8QD1yt8D7kNTaX4LvqobG5e6FuCYD4uavxD8pllL3paCDlOIe0TxmDx/LHdfkS2glT9bfgVgV9
dJRlsrMsvmcaEPAr5pvGITvAQXkd/Avi4FOJ/g5On+3A+aspIDA4mLfKeYGXbfdSMSMkUoLUD+qo
eyvvQKNebH+XdWLryHp8mm/j1spcbGdyMJiL055g1MG1TdWZtWOXnVQdtyc+Y5gRRUFmQXmL6zjG
YtE8nmqGocH9iKLS3TXAtId2YPZhUb5nbf/Swr/vRzOtDgpFjqSeEZYz1mIOIuL+kahCdoQsTrqJ
fODHxCcUf9pgy0JHpY84qr9jdvsOjnDxg5pXkUBiYc/cNVEVHGbpi9cqpHhKV2OP4Q5N0kYs5uPl
rOkPf9VojO3jOQ1gQXRDSdBePLedJHL1S1nD+ajJhDp5u5kwxHO3bP0jolUfYSLmz9gBPJqxXJJ1
9vQDRhQs9kjFg7bTcu78rFSNC698slydT55BpoTWn45/NWdjX/fnFLOWSC4hVr6p3FITm21kaKi+
RJXJt4sSPUjauJT9N8jREQmYueAvCqxHk+SOG/RjMMImVivQgGbzcKF5atUmoQEsS9ViC28i1NiS
D9qOvgyAk8pwD3OZ8sFYfWrGLDpJmMhuncKYLYcynGZH5CE+Ocmm60++fCopv0w/931BQsGZcMJQ
0Y+I1rUrNskMghT/mdqcBnBmc3lvShCtOR+/XiQbOKsyR9wAj2WPhvV44MfnpLqPraooxy50VzI3
cJTSt2QFafduQ6+oK6jRRc8pjPBzKow/AqXJIJaCN/rwe5J3265EccNoANaHa1hUQ/SKenn9yJmk
scv/jPlI16h9NnvNu73RJftPXiaj4VfeZOB7NFccmdZNJovJqGImYz1j1qZykdlSoFBI7fbKbd4Y
yv0A+wreQ9eOTRQAVX++wHPheaK+dvEdeq6oHeNywx2ExVFX5Fmw+LirEz8sKK5TWOTh5g7bAOSW
QnDIqqlQN5iBBKSMYkwUkGny9Av6tdP7ar3NqYCBI2Fx5w0fLlTfPCH2GO/pUixdlrNtgrwas69X
VK3geYuvGFQJsW3/kkt8FEphi1e4GrLPKnXTt6kBzgwF8hZNrskHQoXT9i6FLaAHARj6vMVchZ1M
NMxWS6FEnYAABvbs2SY4wEhA0zKgbfRTbqJ+SqlqNRCLJ8NO6BokG9Qz1z2XWS/I/l77PrS+yChP
W9JmLC8Q13rn3hldfudokplV6xoidRtMl3PzMdp6F3l3ZxKTFjmHDOkx3XN3pXC53iaqXDzipPHL
oTgt5UodMji366SJGzU7S9inIZC90Y50jdwrnT5GFDYwyy9Q/2g9YFvoN46O/I9a2uVtwksfvSdo
2Ktzmmw4PPl64eKeay1QDxlh21SKTE6yuGJdA4XWhDYrYxucxItGM72kDTKmAT05YY62WlQhrCGl
1PSzOSanVI6aXTShhGcUvR3Sj9JtgR7WkOFa10nSPpFi+Z4VNYabkHMviULqnSUJZgxBbj+LhaWQ
x80yxiCXFXHBqUFElnT5YBmCmIt7EskKlDO8U4wbGa+CrPpv6OG2bTBhcH6Bv226LY/OhNku/k5y
95t7uJQ5F8vZPYneXUf4Or0m049QQZhSyUtlnMGfbFlqCGdOA/f+Os5w+PdqQhJf+bk9+BvKwBy7
wSVWG6V3camEUsn5nsj2wGJFd9ruoWuDNK7ZSXQboQ8aPJ4brP/ktRnLH2BwCZSfloiXq5nqJAJn
/Am+WDWh95a7VaOqDBzHEP39Ji1ebMGvmAodiGu52XyOg1U/ME8fKUTas1U66av3CekJWrN8ykq/
wl75OSDD+6h/dH5nse2fQXK550w/ZYyGQD+6j1rsh6P8aFNDEZwl+8ZqzX4UeRdsEC7bql8IYry/
NdRIParapxaWYChgb661wwHj0jotTvL9CSlPCa2tfGbNng9zB7kxz4Or7LWFwQ9Yel0qW+W6bvX6
GFLHt41KsMvPUjHS+VFhLbY1X7LEt3Iq6aCwQ47CPfTx5rZKQr7Bfa1kSxhVjeVghpvswNSrHLgR
4WggMDntcH0+OEa/6Cw6E+hdFUvOQ6ILE4EHmoAUkJX9/yCVl5zTXnKNPpLXT86xhWRuV+u71Vdv
An6JfX2Atc3fKZaxNE7WIi4DsS8nJkOnc5DDK7yfh8Pl4DeLrlOLjJ9K9QhUFKa0iFY6Yjl4xQXN
UaRUCHtVYpGZypmARrCPF935uqQjsy6h7Y02sR1MVgp3OaWoqyn2N0PifwkCDgUSf2wtd6aaRMq3
yGhSLOzBG6mu/depT2FfkIyueU+3kB1vn1m/68u0Aq+Q1pQ5YhrHHDMx2DZSGaoHz247JUZBV5Bk
7TCVsjFViiTsKS4lj/9TNzsGblNVNgbf32VcMdlUMxZD33pcTFea6XdQs1/H00WphAGBkj5o34yw
goBHZrxGfhKYkL3ojWW6MB8/KEN7ekW6ZDQHznJxMytfqw+aUFwg6Z5GiPqn/ahM9Crx7LV8swDk
G6zTZWYAtitcFkBDuNqKdjxy6Rh0q6aW4Qkb9/XkSHt0wNDgPvw3fBLz9jZu9vsG8icaEixJPoSu
q+w+uSMErgyUMCBNrHkrmUMxjExS+Gpl2QfR4MrS0J/e6GUtjoWoD9jktiiKAaLaLAOo1Q1d98zj
NiF5X4Q7Ll+zo7oV9hxn4jrCGY7mzEL0RlUwpkrbISaMg6HExScNZn9ybyh5N0PbQ09UF7Tl0OkR
Jkf1v5aMpnvQz2A/Rn0+L1L9Yq7oN6/NWIjBD6mqXIgTZtrTpZ6nqRCwqt+VXvehhXDVrMgvCNEf
hOv/ajawmtzWGdmGbVOgzTJtWTpK0S4UAXjBAS5yyh0nIeYoWa7lASWYmnaBinEUE0EH5RgOAsmr
hA8R7Zb8sjQcjWqYmgJiiK+fS4lMZj9+o6ZsYRV7tZIaRQrmwPFyYW1ey0YmQVKzrCoEGVSCIsqN
Bl1aAG2LXizNXPOEAVsFFSe8ZwHqRvGdWLP8/YXFC+A5xQExjBqdSapfbxFO5uuGqwK0WuNsAk3O
UXclc7LatJovIBXbTU5bkBZAwgY6jlg8x4B82UUerqtKpQnWjXbg7C2lAhf3g9jNriyud4D9CBod
sJrkH8UioCZdaIL2g+dVmMqfMeUAzTJ2NpwWIeJv32XyTypUPlIhmXCBOMNWlBnjdUgoJ/TOEm3h
JbJHRVlVEPIMMis7qchn0+PGi7jBMToMTr9cIB3Zy/D+ImbJA8v787wsOEF5i8PTYhna0fIdM21r
XlhYp98Jk2lvo9PcFcW/G7uT2QPpd5H+roSngiTBsYRlT8E+Ki98187gG9WE074G1SQpp0s0GV1e
rek2jNy9oJrdR2h8DpDUUh0nabZEMANRL4GLbQ6e4P3cV7ekZrQFCknRJn90cmorE8+D+BnB13IF
2x9OyKRJ/H2cghTwqegK3qfqBLQy0mxhqTdutUkeoBhzeaQApyrlM0iD4sR5SBuTm/l6HUoDvniT
byeTEbLsuWq9osJSSlrZvbgxl9jMnB/p0kN/FPwaHst4yThV4juINQa7GE59fVAcA6qp4vkxivnL
Ed5fK+4fAxbNG2/hTikDo4ORrh5NnSHmUEfLxlCylF+5eo3Z1YwjKwQrBWaLG55D8zasDuD+xYz8
G4KQKYYtr/L5c7U6eJiJLfPCguWwn6p1mXM49pbumM64i9sO7feSYt0yzJexHHOoS9kmrQ3jXVmT
WNOedf6TLRPcDYnXWWi+53NwQwrInDTavk6arxrd3T0exPCQ8dIE2iSzqpxDDoEEdfbViyu2Myxs
kuHV/j8a2eZJL8s4wtjU+70yWQaR6Ncxnag39M6uw83tdhoKslVhhhcbNfl18feP/8S+LvjAcHUz
w5UCHAz2l7+5AndHQGvuocGcNnVA+k5grg7xH9y02cpZkWDXdvYxV4DONa0vho724/cp/ZY/vyWB
1LWKLUXq4zH8KHtwixokpMB5w+RPhOfzjtrd3sPIFJwABooltr4Jea5TfDDH6uNQXinNhOzeVjAj
2mEMp6ADQewWE720iicPuaBBkvjQ9f6tLn0SyfJPx/FjZFpt74GpgfrxhoVO2Q4QvMOblJfB9duk
oNVT61tbv0tGdQG3ItdLP99FMzUw2TgaIXoE81LuHO8PhBhBYC/ZdQQGw6F2anR7DbNy/TaFeoDW
t+NljV9eRSlgd56On9F6PVf6mAzuY81fzX7REovp5ZSjA3wmUZ9SEx25f1y4UYjFMmviYghmSPzf
NktlkSwC3idVJ+9/Cx8heuCjNJxTakhkqUbl8n0ONdgV03GbzAnjbHgIEDaKSTbiAr3TLLOXq+dN
jh47LNZ04DSs5EgcFSghDNslg7ylqZHazwYlcmryEuXMXkUfr2S4zmosflNojsEgKUKXd68NgM3g
YDBlUhtCjamvmgTUj3YD13sOvZVTGD4vRLibhmpQeeIZTnDnSZQK1T7N2PskwxblgYumGhNB2uJ6
F0Q+LIhtgk0dGRI8BvZ4ZneAsL2hqq/h/w3gVBnVcqSYu3XsYqBeqxeBZolXU9noshwY5EnJHtCh
4LbOGQ18YHOlUa44gI+cuDqk2LQOUSvyRfa27Mw8NZtEtGFK3J2+Xf4Vby7+OXEk+Mj8lKiMfLJZ
5/bmxejmPjzIbI1UlNqpgu4eMmo8wDNAq8JK1mX2eeJEOBU+SIMn9EnGzZBdCs7gzpNJF5AXcwJA
P9RQ8+6uYfOAwha+uXamYr5p6uz20UyQB90YaGLXND3MJ6wdJ4omhz3ZJpEfzk7kTl/Xg/uLHWtw
badydI4oRjAV5tCaNInXrLKsXyD8tkunIN8YTXoUCPp9PUcO/e6Aur/8V2JdyatGzYU16c+wfPl1
138JVJojG6tDvjnag4SG0nV/prG5mrGRPK2Dss1UxKkySi+pDwETn/zuizUoQEEGBEtoYDW4PJD+
y+HmMePE4CUCRCl/oh/MNgpNaNute9xdSkQg+lmBMgsDudifnCY8gsPhjtpnUcxLNK59kvPNaU5C
PVQ4mzZABJVgP6uNXXPWLmaY88BV1nlh89wloeaF3S2mBYQJf1XOL8g1r0j1WfzFPCycSm5nTfM7
JGZ3/TOTF1Cf91TEcFTQXs85qsF54INodetl0P5EovRrPLo8CM5nLUP0BFXsrmmhsw1KbwmJabId
qcw4Z1ZGoIuY8Ln3GpyUuvFLFA0y1PNLEUGnFMvoc2KWZUKTFcuIKmIWJ32cKrJ9LyOIwn5Y5j87
eCen5rJ9DBqrwJ0qmqv9A7hMtd8klLqPkbkcFzCxRGhZtwAHkxVY/2Yohh5OykH9h1oN5K0XYrG0
g5wNdoM8xnj5RZPTGR6bN5pxWtwCZAI5gSES+mZntqwJoinYhcW8xr0nGoJdzF0Cqku8jiSikjYw
7Dn84OZ7HEubd5X8XdOj57LZekdu23HUATi8VwdIybIMIsRzmdcrQuiWRwHLtbQ3rC9euYQABh94
z0ZXyVmoxhe1Yl6jckyAOWYH9Wc1xEskbaFU/F9DHtsULCFsFRfygRv3HnxLhRRpZ1+q2r3sqfL3
KMlmip2kK4nVrEZrqtqFxXeN94ljJtTWbETEQ/InoLRzQM8ji/CuEcvloDYiPUsDVsHtHW+ipsZv
GBO0yi0dGpy/N7eQGXOdl3vu9iK8w5PaTS0hRgDJb/ArHG6MmvU7cZdlyckDfghOoSdvOz/LWamv
YhHn51BKup3b/Q3MqojwUxTLAVr/gbvNk8ne1gcB0CWqgVuVFnN4KnpFtAbZ6v9TDk0eqJq4LOb+
H5w6fq2bdueZ06rFKrjGhthswBt5MawpoRuWT0jPwZGUZgsiCJ1FzDLxIEdI/PZ/LkzqnNBZXOr3
O3+bjT162Ubh5O4kYBJknma66WPkrtdNcmGweTG0zdvGGy/ahay8DmngUki7Ydze/BYgRDI8gEVl
Yn1Fk17kG6fV3z8igHUuFX/90ofi5yZt3rwPsrTXkwflaHDBUKpjOZPfqBeS5HXxpBTcnVBo4BsF
O3BeSBMENoKvRyFGAbqPUrrWZLdG1W34enSR4umKh8Q/0hyU3tpKDTL1XMlUf5yeybyLVfY+ZU/D
CtXS7KfOVquNvh9pzfHTctCb1PkZWasJDEbLpU4oFCiZ4mkdWfax9T9w5c2vkND8fKGPKXZQpOgX
wBxsLNU3v9z/Xe/FH/7Re9fuC1fc9NATGGUzWcKpt7O0b7KWBvihyPA9A9tB8FW5EXayKDXie3Xs
j6GgaAMTghpM20sjU5/biqcYUoOI3WG2Ea2Oy1dGX1ALQ7J0L6+fDz/WCI4e5LsO1AtpRht7eva0
uZeWtfvrpnzrefHxqJ/xb8XkFyAD9/wk/KDt4/6DSoRtQOnL/jkocJYkDa6mdTEodvG+bTYiyhYb
CT3d/YGOfeoLmDU8vq9DoUCHrPi6P6Cp/AGnaeVnlg2Hf4XQ0AUsB4Q0w9tkEwrS8KxfkroE0X2+
ZOHr2REOzqSIENloY1aicRdhjPpcWt8Lm/QddEWGoQ9YeG5hldp0URvDnfEiKPSngDHQ3uldFZaW
MGEhqBXKi1I4FZcTQYvGxWzcNmIE9liCMFvUUad4ZIIJ0jiFbORNWeeSrbwq6vPd5WQiHIUmCnvf
MVBH29wj/YFgde7fAkFmSEi0MMX5qKO3/sm8mRqRm/zg5cyZ87oniD6wBlaYH1GUXOQPqn18cm4j
u6gLF/6LpHFBEopTwdHRZJGF0TN18vV2E4/Q2kk/VyxrSsfsCZnT4BIttYwVrKfDuNZJvALKG1QZ
4LOGBAOfuozi2nmNPd9MqPDgjqrW8umCWBOAysgDeCSb5oR9JFPyLR9SFYuVOVYj8PjlesYa35qV
syYdbmouuTgqVLCzWRTMJ5Re0DWpAzxLdkg8ax/gzmSfW4B4f7cWcc5osm/NywoRqGH3a+7B+476
hq+13innU7QNP0Y26GJGvsEzeAXdh47tHcVLfvrzoKeysM22/7tEQ2s1+qHzEk28c4nWJrBRKpsO
hMapbrzAub1+uP5lCz8liWgcHKJxfwswGTmar7ZSBQAdslUXPNwHDIUW46fIzAiS69RcFoa+MsfJ
SGKK6seAepZYaLBuG1WOiFrPIM1SQlOH9i0gFSEl/Gw8VIPtGj8SLMzbhSnx3giP7mjurHchUJTi
iIZooc4170GgtAIg8qPpY4ga94iQUBNNgH2vMdmxNaUN4xE5Nr5fQXBNTZ5GhcgO00rSLoqoSAsY
b3bjg4J5dDl2kx2WpPdvBQXQSkiRbNksc6UrJ+3teiPc73xfdSD4tmrXG37qRlMyDX7U0/VXdoea
opFOkpWiYRj0myISTkvzRMNrLsxraldw8QC7j3IuAsyJKGOhUaN0lwZJzgLX8p/WiTRVU6iwZWKU
BwU5aRmdoAmRghTA7tuX3fNghoKb6eq1XhaGzPNondyMykk4H2QMTmoY5jlTWMijh6DpGVucV+YY
0RqA8rGn3MoaYOJPC/ND+m1ukpvDw813ZLOAeeZg5jeUcBeB0tiABuyKKo1wTzbJ3lk0asLzQTJ3
Eu+VoIBrvfE2i82TS/pK3h+ryzJYqIbkYKs39T8QQh5TZ4Cu5it/1dE3jxlB35wqaZzNC1yrtOK3
o3rJttl0NJFZrD1ORqDrr4ygHIC9IF8/FT9MFUmCGZ1B4Zwry53l+mFmMIz67mj56y3ZVvuc7oDs
XFGPtAJ3g86gKi+jkHphxos0rmEWtOmAtV2pyIVtetNz76h9fDDgIpGLV5HpKU7Dgcdp8a1HF3gs
xTte+gSkBwzRSr6OsnJnpFmkhei8s5lPH1vrFg7oTgPns+2WUY3x4LteAcvlAk0xs3By2YfrwDg4
tpSWMEowMLmmZ7Ncvz5nDMpACEkfTpC6ohRS0y6KFRpaqxDu1xi91W/frvGUFxgPgj3A48Ag+Gig
vG6I6lXFZkLFnTbrvjLY7bZMDPvVF2c4wwn/sLeKFmoclQyiE0fLG590sRQxAF2Rtqxhis/sFBu5
1pQhbZ/1QNKx7wciKIQVJLitPf0B457U0jyEfyA9DPA0jRneVSWNJzEhr05GglwV8qEuZI3e1+2d
NZJLBwfgJ2BEAqPu0rAHr/eRc+YTHGCSSGqmWjlYt4+zndDWwxF2dl3XaycVnoQBoR64bplmH6SC
2lX94I5ZSpQGM4B3owu6hzCcnBDZICL4tfvKK0qUNSghAcy3zojKyAiW+ngA9LoY07R39dTzq+yM
t5PRobueh86YVt9Jt/lPwRE1OPTCApYSRFE9sf4yN/vVxemptn2aSyazBomGloKWl13+NzKkEZgn
nUKMGvzoOlXCiSc0y0JSEPLuqdadpPW/WlGRWU1vNa3kYWT06Jy9dun/w5yxuG1w76fgWBndxLMQ
LypOjGP6UmKE4SZfcbagCjISX57ZCQq3HfqPlB3PuR8ecwjNK4fxD5xZ+3+QNY+AuVpd1xf+JVZf
H2vDFGT8Prrvb6SqkucHD6VVTe8sAoyjweN9CtMZ923poaLTig2rUjHNVdxNosjZYDFZkT26YBdN
lEkl0v445Pi+PDx/xe1Re3o38n14BtmHYrileHYXiWr741kLNiFpPmt69m3MEwD+gPiEdlC1gs+j
FxjDBgV1U29LiXQOJ1XYA5r9exutdlJ4uSXxh0/6Bil+kAy24O/xNo2dKJnd574F4vDUgnvyz5j0
TH4008gQ7UH0yaKxhniva2oN2L+tH1Cq7Z2kFOqadjA1WLhtdSyQF4/JkHm62jSCL186GoYbBU1i
PF1f6meR1nTEeUvaN57BlSGFySfXYUGM92lav/kfTtTMRM2TJPvp8MGhvG5EQ9Lji9Tz2jX8Ig4h
6euIV5gvdOdGNIh2xXaIjZSPAZSW+ELUZlgHKmp6Yc7jxeKdDsLAxuFS2nb/l/L5sTCE85FrOqA9
L5hUXl98OfL6mTCsGKGn1stRpeqL9r+bzPeSWJjkrZnxzheEN5c8jWlmlQnQRN6Uw9jHaLgGOGJa
Vy6/BrswWY3+pVh2jaHgIw4tabOnZyU+zDOHSIX2CCwCAzkitCahSk1O01G1CgRhznr9U73X6mFf
BimO/GXUPhzcUpDIz4THBsXone+p+9ErNtvhBqiV5tgCBO/NCsETSG+G2dyyzQgco97XdScn5vhU
xcmHsUPwS0j7EnSDwQfrmnlmbnocfoM8y6d30kLBQIGv4VVIqnIGGi1j4vgVrzAGZeqPjEsEu8TR
YeGOStqUkz+gADpSwFRz4Tf0en0em9bV/fM0q7aJoh4g3Rhmc0y8T0axD+In6GlJroLnwe0wOcLk
KUssuBkYEYwXc+a+iukTw2ODLrGjjWArA75DZqEXsbnkJRk1nHqsCEyG9DA13oeo/jsC8DiEnAYd
d0/+wJJN4EaQTW9o8R8noHWGfGngeW2nZthpaJfU+7UuYA2gqGXmrAq/gFYKIqYsISR9dczFNCT6
yW0RdVnRlQGCDi3z/CDHoqP6r/nDPs2zl9ptnMnCf2SGdz7bRZLWZ4NuUGDpGGRR+envA1zAF7Zu
CyqIVIqPKhqEJZSMwrF2ACe3IMYMPaILzL0lpYd1mL93yWA4WcdzlkWmf92Kv0TKMf1ZhfGGhpKv
EwWR43RxJYaZqXt7qRhfLSYsCWdzoA+EBcpViXtr6sttr7PzH0wuTCkHPGi8orgIVqj1MtzsJ0ob
Glk4PYo9vsW9HduGYXs2qNJs/1j4gA2XtwQ4H07ftnb069ElUbyvWmUEtPSBS4LkWn9OnbZ7P6Kt
/MiHNgimah00DjN3cQe97fEWqQYLLkU16X6OSsck0Ef+Aw2wsn1CrI4xdPu1y/884kLiUtf7dFI6
Femhe8Q/ohz3yNY6JdZmAdZgHAlFSd1nnYZGQqLCEGPGIUJ/8lPIvWhB+InW0sXj72zHQjnzalN5
WIvote8mM7zPNwTt6r8KMN0NeScp11Yg2cYviv9FkkNAaCcS4poVzfZVbsPacdbenf1iucT1o/6l
m2uEac9Fbzx2ljAwpRq6jK5BEX23tj9yCRlIwXPgQefzR1WYDBhBfHBeEIc5q7BA7m8P70tlzhxG
voB2maZOgc7nTbDSkO/ssr95BuAiSwSKFchqbu1XsV3hf4xcUsuaFMjjknxaa+Ctp/quj4ziTOG3
uk+Z+apCqHYmArOTbder+vwmlCgUypSuFGbt343xs8IxcH48U8Oo+CtHZZ9HovUUYMd/l1Ed3woS
Q4YGpqrSdm0P3XBr73i9n2NSK9UCRlyrkd/UGg5ZOwc90HT1PuSc3QG3f6bJhyOKp2dscxxyXxfT
/Ro1fIfVmYtgo/87D3yorsXMusthr0EGMwKihSHVcS2YsubvnU4tRNxYRJ0ym9qsdnrNIZLUhQdB
t92dtKGJ0UlB0F7tms/+f8H0Z7QyfprWm67HGUc1GgYcysmC5aL1jiTG/jOQt9fm54MtRpCSJ0v6
iRqFXNi2v58TPkefyd14H3kWke2l1fLbKbq7XuonB2AfuIsS6/aV8ViEyp848H6tWPOT5kgNbBkl
UGnFIfnu9LfmlP5BWTh+UQpba6XbcS5StFANeR+RZJEnhwgR+1XBC34cwuKaafzKC2Stl2Hpm2jh
W/ackmWYLHptECxPuiDw2pBZTxqZQtK1z3nADDLfYnLJI+vP8XTAgAxYXCozYGyFmdKu6Smeuv+W
hQmghHHC9GSRV0NpeDHWvDV/v6sVchlf088p0+LUS+rECiwfUqh9dNIn0Y28eepp6Id4rMdOgPuM
rDxJsJHa2/rPRzvDfAWrQagpOC/Gi3aAd5+m4XEP/biaK4V0PKSK/ovt1fKfuo/dkwy5HTcZdyaX
RhvSZafvFT9dJPZYJMg2nlfe24tLlFuP9YoBZo5h1Zd6jZUHrVpYQSot20ZcUyvuvrJSSqY5qqcd
eNvZjZpP7StrfURCLJ2oTxcouEKM8mD7oAD2vwisvaAoPESXUwotlwcFOgMTllluAqfIlmrWRNkr
k2aPlOmV0DHqBCjrcupJ/x7UjmVycjih2VF13Rpv+aekDvY3erdfBJARNCTR10+8JmS873Did8Uw
0v6Ql+vqPi0nJAhqB+t6igEjb0gT0tQjKHILVyKIN0WzHXoqKmTdb4fnrgjHywLxJCCSeaTQHJM1
JOtCYmcsnsJ1qbe8MNP5IkhOuOCybd/U+f7177tiIG6HRb/pe9BomjskMad9U/c2ZU33MUynrz7i
AsrkaEZOmJhHWe9Jj1VwJ312p61B2E57sJuaSke77A9L/6+7Lg+W77kB+QHEL6+/00V+h403mbCp
685U6Fay0+fefLrwVUaHWymX8Vppbqg5KaG6VZknaSWv/3YeSCZZjzDQQ2DhpzdtOtw8LjnRB5iP
W2a1lTTTapG2KrVu83zN0nHvNylbDj4ZJ5wP+WX1qBIedZokZF/8iz8Br/cxX8ppTSiom8e7OFeU
vkf4PlNRilqaZDLm6g24GIQ7nvb8A6iXW38ISx4MiVMRe5Y3xs2Ht1yZAWhujaNZWNRYniXLV3fv
1aPiQULeY72M7G0byIoyHL62TTQGeYZ2ruwaj7GS6R1vlLyEu5MgkUczPstngyuE/q3nFuulO2al
deSq/Zp4AhDXSRGojxtubcR8gUkpSk7BxwyC4QJZRJb+r/PbMU8BIGU3Q2YBatdSlh8G/5Y9wxE2
iWeuciBpbcpUwffr+CCAMjQepcrNk5PIRPwAXzYEOeCo10CwbeNnmK+ITWwC14HjfiMxsUY/2K0J
ed5ng03r9+g/1eQ+TREavnofIUd88dkv+3LBP5pLA4NbFT/aqgwB2XQBFk7z7NcYj0G8SCVELlWT
BpNy+6ySsDdLRw/kII85bg9D0fRKplFhW3dX1zdHsWyk/fpziIzbkrLICDbvdLi2Gz+uobg6XNni
ozrGgnq4F4oZ9ayR0OMR9dFl+y5qdDqWxWkjATOsOCKJ9KE4EqkrQQV2FiizkpyvGkXJnYxTfCC/
R4d6C8nt60T7Drbj+PLxX0ujyGCOIZnWlfWAKu2uhQmD6rNpGOWoYG3UBUqYIZA/Yv4aCTM9Cg+A
sAKxB/auNzzDJCX5z4l9jnD7NKxNU46JxEr+eYDwW0CJbdP/ogDezoSO0NlBj7zdj0+NF9Y/ovD3
SFFC8BJYIK7NFs3WTPrn4Ir3M+wofgLJGIEj6/XnNwInxu3zrQJBK4Gow56hbZ7kVituNq2Jxg/2
xrTIv+JeJVr182xeryhgx0knv/M1iYXDgPo/ZJYONUzuc+pbnSKDbxizAzhgk8vJUI3137qPEbWJ
V3m0AfLN8WTu8no3zmMG10UudOzNvnbR9RX5dwS20jsIsd+2OqE4Ey74DsP5XPKWeqPx6t2Kldln
KL/VJL3wDtdqIK7nZ7eNMBx5n65a42zklVqyp3VwlNtpSzt8PEMxE49IZqMxuVJgR+CY9Yh0HyN+
jkfh6BZAshQZj3pDdhz7vr9qvwD8GLTeEcyfc5CJ91RHQ769jQY05gqsAxCv22e67+kwvVhOCMha
mUUCCgztlr2WfehdpaYMfDC5I9B/aBtSiLV7BOt/1j8DmC8gyp+7KSOnfPkjo40fODNEkAHajyHS
yx+WEpgxydQhM4e97JFPWjya3m1Ln07oRkhV3PDNvIgrsXrsHK6KNtwKRMRpYARPUI1Ki4JzkSu3
PLzmgQeQBm6ug7qTLpXEU1fz/jeUAKX6ZyzRdkVttvs9pHkoQ9DcU+LA6B76HlHxHk6kgIJ+/dCP
RCL7L/ZmMZpFZq1rbmzfbwqa6UAnQNLxuA9VvWCrB3DmJ/sKIVwtx7+EPcMsyR2VCqA0tjq0bJUc
ox17gv39Lk+m0ojZV0QrD49horTDJFKAAusje3lObmi9TxbySr+7cAXqBpv+S0LBSA3CaFeRc1yl
D1nALfMcUBXgfhPtCmunqqOkGJjtytNlk0IQQLDKW072tNqngJaEsFwQ19gaugHHW/eiErlVEQAg
ZvePzpdNXErYEuzSLB0Wn5CvsTmoM3EkqkkaYSYLuX9FYFqIlbxBY2VXOZziBbJyC0q3I1TU9f+4
2MqKV01R9byhxUnq60bxedJs42mw/CWTsolAJsoUfWOshqdUBadOWwMfH0TmFJ+Fu2gSNsr8St/p
CWOniKi8MS5SqEfRxFzBMwZALqzK5qbxuxXJYAusE8KVMa26RQYrk9jQZES0NLxm9bsXqeEbnBlV
9RcnsUU8JcKvbgZn+bLXHN0RiLUkDuSn7qShH293j4FtBT6MWBOtD69foDFvURSykwnSEero4qKt
S0AVK7f9i8CN0PG/sRPg4mipjuNzs1+acyevQQGMn9hxl9lSjoNKHOA0x2qVPMN5J/hLf48f5axD
NSuWOdgjcGlnKfUVy13v8d++pmEaoaLpKTyA0zWNa25vYO7c5iYkDqYlUOxDN31Uqvsf+v4reUZO
tp2+AhDo6h/uWv5uJxyTIIjQwZtrjeAMwWGkNhupa7P/I/sg19RiXH6BfFvju+dN3OdcMYJXlHdN
HKb+A3SaH0xyqXKD8GJGQV95SNnr2tG4YvR5yztSGq+G2SYTgzk3XdK446qZabOEReY7E4hlJhFM
EU7NRg+KjOHaWtGMJ3hy4AeIpzDGN4uLFfUcn0mRYVco2m3NNITs+MVAZk+rR6kXRTNDXt8pH5gr
+mRU3t4A2ZpAWWXxnBwkLMp8I2igFSXX5n1qEBisloGf6Gcs1E0eVXuQavh4KGinj95QlzSNkolN
S11/O+h3ReSmeRvUC+1CmIGS9Xbl5ymbe0EiVOObK1onusW3KnvE84lpxm4vroxtXm48Vd6MQJnf
SBVaSfBb5d9VcRwTjmn7vbdnAcz8NGHt21bYXb43b780r/QDO/E3KsbIibErX3MrLEeFG0pNIbJq
TqCjYJtXXgwcxClqSyWDYteu7irLKUohrpaiND41PrywarHi8PjOzjig1sU3A0jRH/HR//WMJ1uD
kqwGEyonUL5dahU3m9XytrG38/KYpXXobvU7CD0GuNPfodp8PBYkP/zNbT1HZ5vOWIDuoAllXear
c8dVs0lmpwLGkVo2jDZxarArhuJCW0U4YuMmPHAl8EBkzFJWUpY/gVXnLmAm+iCPD0+asBS/V7pp
EOAz5G0p35SICUjs1d3sA2PTYEsP1Ums53yqYFOtuDZVRujnstXwYu3rn38BBL41NFK37r6yN6g4
o7LljMm9FtjdbRdNhzqHpHKTZq782yMw6yqsDPbsOvgBVfLn5vA24PQUwWBsEKxScgMGf13ycJHV
Ngz31iI3iuvV2Gr1OaiyZUjlrywTRsCDvSkrcw3v0UCKZ3xlRWDBVcL+i+eA0QSqUa+F1yrHBcza
QbGOT8G73D5DMqcv0n2F3PcRC31JGaUBIRK9IwIAGbd/wsrANFbqnHyR+5g2YrqEBhNo3ZZCUp2D
RN4GNhgcYkAgx7eFGCy4fpOG5WRuPc3Tw7AivNIkZ7eRBaNO/aPKGwc9UP043rWTxFUJ4fpUjTCi
hX/eL05O8O7rfcP2YykL7oA4Z6/IPNvLMz5mxXhP9ofO9HHcCnUdiTA7hhIhWa7mewhQJi8lyg5E
wpgtW7yowQ+GqzS2mzfrDTaEjaywL2jCk8jsgGcdrO+FJfqDW5DEucrUlrAw8SvgXT+0scF6GOts
h9W5SoZY/LLAtQQedTOPG8wN2zgdcqB+1a2pZzVMK+04td2Sy5/zWbeeJ56r3aegUT9OcBSiA5Hm
IvOgxxru3K7W5bdRHRKGXyAr0YWpClnmnNBByNlMeu4Y+smN4AAOSzXJnHbTv9m7umEZDl9BNj32
Dod+jPmHOahUBpbEbG93pPVHtHUgeDSQM4eAvEYG6HABO6T3CUpck3PxaqVmVVU7QDYfQzN47fc7
dDYakI7HC1zhJhXiHpYQBQDOo7vYaVI8IpodaZvUhG3OZ7943vb8ps8KrS6Iaw6Bf1e4eO0RQMaQ
tfcH3BDBDJ3aYP4ceyRdhEYKa0e7ebX9YmUysiEEZy0y5uZK2SJ5IGYPNNUQjcXeoYZ5S5yuHqiz
C4EuUGXFKmxNdOdnz7NfOZkShBdgjUEzZPM7DgDg7zYW+7c9zN2KIyTHla++lv1F7EfdxeXFTUhz
//e6H9DNfJZIwWEzFnv1CZ5R9hvXwQgXBPGjRuauzT5BWZUiSD2CYaxVibUtan2D0zOZNJB9JMhy
a+P8+aSU08TPctMuDwk7JXeTk8QhVxrxG5i6urgi0CyzoGtuLG1QWoZwKylsqpqvdr8O/g8hcgCH
ih1c+U6y49cH1IW8VqRP5HFGf8aSWNOtr8Yuzv6BK8m/BX9EzEtlGQJWH+AtsWZme3MfQrQCoxyU
G1p+E7xQzI3OSmowYJl7BpPLMN+gpYaxoDrT2lvBTJwk7o7lZGeyF3H3JOh6NW5/ed63W8U9LE08
v4ixmNYKW4hpwTX1h8eYgc9bvXc1gk78pCUWN5SqpiVdIL8OlWl6s0vHwIAuad7YlVZo+SBwqHtQ
Hc6vkyb50Kul/VQluHMVUYjBAidRjwvsTyBUaZLNMjP5iBneb8Hr04nr2oRJQtvuoMTZenMAP9yt
quRL2sGW8wqVJmzHhSHb/ao56e9gZd8g1/FPPbCnluI5ZMKbtklw6lDZmNcZxO3I5RlSP0ZlvRn0
3TqEwBd1XrbcTXGG5zV3X3l1K+tlyDr5yh+D+llaXLVXuIADvgo6CtJ0BvuBQMeyvEiULdUtdtH6
ex0cTdsY/Dq6K6nNBUKylwS/3Yk9/6NF8C1jg35UUg3Nz8BB02TDlqL34BpEVSUbC4uehgSOa5yT
qZ0F75iE7HKTU0CI2//lnC0Rgv96DGwyYM5tAGTDTKcxuwYHJftCNe6wNnbcUiPWjeZB0u9RxWuo
l0bVVgZ7wssp9COu3LPUrFWr9qiX8Tm4ZaQVDw1AHM68BRHFq3eJvAC0IV6ihgjxO4DGNgbBPL/e
QhwbnF2aGB2JKremRtRctMm1j8us+chKyK9pj1E6Po1u0UJ4e1JToOPcLQ2u2pbygQLKn9qw/uwO
jXwcFgoHD9XPcxd3q0FPQJd3g9Twqm3QVQ1sjUyVN1E/IqrOuQDHdJdpLiV7C9IdQo+Sjm+e04cr
7jO/GpvOC2pYK+V/wq+zeemEStAsyTfOHek1Iagh70kU2IpI0dlpkaMFY8fe7Csw9TNwUO/bpvWQ
wLNAqrPubrratZ1kKVxb4yZvYXV7RiilGweoPfF9f1J2KaXEkBtz6XxXORyb3n1XWGfX8jlQ+yIs
GVOIIxPwEDqGCTDzxRag9dMZ24T2hR9KYXiJKKCQ4foTWY+6m7aq5EqYNwSVYsFLaULYNb0Zooea
ipnonN50ImteOUqJXGry2W4o1MPNYrrReunZI4A7fPfm7yv3UE148azMU0q/gGxh39suLT5QBEkt
OxcscTaPt3y6wW/fxK3YrpInWzT8AsMxWolBC6/bnS/Xj7AeMqwr5q7Y9ZoszMZ41guKlXNevetY
HXDeniegH6QQiqTIzYNDdSRr9yOinbpMI3K4WA7ThPpEHG+rM9MLGr+EYbbCjmDmWTVUHGKI+7bJ
tX1xAkokab+f0kaH6ug3I7IY9aBmQrFg+/HCVYX288+hlL4keIJjDOoP0mFZtv6iM6JGRFaqPKLy
7GTHELvH7Qa+xmxgwzKs6jQKiaU/lENKGkP5J5AmvPiju7bDn3rk7YxO1JMuy+uRmG1uITm7bJtO
HpTQU96z+Cc+jibJQndTkGLnVbNZ6Sr5NXSQpFaHCL0jzSQAHZGutMkSxkANVgoOcjGQ5WerLrfK
Y2uUMU6hbnZ7MJ+uRNgAiLqL4YJ5gTpMzfuoO/7y2p/cI/jOAmsEmF/76Nvf8P0FC40y5BUTOU1U
2umWu6+iD5VBdoTEfQalPT0RG66HirpkwNUlJ8/LtIMl+xYXppDIcOV+bwr4shUO+cH7ioZnfDOz
NdfUG7bKyg5TYVbTWw8cY/8eb0cnNDdsPKHV4TS6OaWVHkozBKPvo8xZ3r8mNOidNL3XJ1HRKF/q
/mnyoTpYOTWUVodEbN3yhakaoCN6rr0Z/AlXQMjnh+1eNEwNLaezFvGthBu1ra+7+T3+J88egeDa
kXDqObjOmVRYVWj3etjvqPksjwRsO2AcfByVDUi+OffSdJPcAVKHziESBxN8H5nIupUUpG03wwVQ
6Rv1i/lHchtjj7uyCUDDAKjurAR6MO1sXBRHqIN9nD7qBHMqiok17w34vrURoJxbEx1is1ZpCSJi
wbbYbfaXpNZzq+L0hWaJH0LjVfq8xcCDZDy1Ucl0jpBEj43FxFF0wJprXcZqxmj2M8GWzpQ9gKtV
O63GFbcd60/IbGHJSPYvAfJH4jcR711UhXwtTg+0N8RzkN64k7ty08VxeNTQi0hfszEI/VDe2zy8
RWeXol2pCdv6+KIRZMMaeF8FhpC78/gRKDwhWhx9t2CV5p5Ii4O4ZU9OgOOGq5M3/sNlHFVfi7Ip
g9ZjpizBeZkhEbuk6HPKQw1iYgVcaT40rROFfBSOFNj5DnkdBwO9+h3J+cFsvq8V9rp2KyezjYF1
E4WDUg5uLnN0QJGXOwg9BcE79M4vZ/HOl9+pBRJzfr6RzR7IaqcAOcDMgF+oxmB8g2ceS6Y8MdLh
A5/IsEwNp2HX7FaaBG5uvqLixH2VgKNVnw4OD3CfORVgCYD04ThP5dZ+0rkHs+5XM54Dl65vev17
jc8aMZSdq1Ckg2QoTW4Yr1nMujW2nD8zOJABV0AsJZ0P3Ce5r6AE7tycVIGGXvKr3trNYxWcrtA5
Q9T8NhkWOAr01AN65o2PljEz3MO0Yjn1eYKHoKcqQpEnTcTMu05nKTEPO7ixeZzsupi1gcYlMV8p
1UWY2/7zmDFT9ctCS+Rb1hS2Dydw2oT5u1/QqG1G7QkPRFPB5cV3sVemi/Pwds+hqeT5/jLFqZPD
NJiMbFaq0pP9CZVWp/oNvsqW620LTirKxMM+OIZ0acRt9W0Lfvf9UVuZ7ogAVpJzX41Fp/uG3+qO
oSfoLcTnnrwMPdF2oXawSpXIBvq9p+KGmoT5onp70xEtsPPayL5MNMP4JEMTBc3TjQ9EzmSa43vH
qN/Uad2w7XxHstdoImSZnGNkmFfkEAusKT253ypBDyS5XXpZoiWsLDkCyA7qKE6KfoO0z3v9xiCt
WEk64oCYpaVL+1wkWh4XgsOZoIDuyUpqgx22h1oLXLjqKxkd1ktoJY+T8ysD7+heXex8cPN8bP9z
JutqrG51PLKXXfnpAWlSO9AzKZOrw6l00rFGd1FNwXqnIB3FaEFv9uN6cdL6Dvxwx2efxcwj8ABG
GijecYjms3vxI9ARpILfPsVVmhe1p7Ul3Z4VQhxG8kx4HkxNiKfqtTzLsOH0fZZZ4vbuPtH/aKWZ
AErho646Z5NMKkN++b/7Ndh3bg7y/rRlqCfXmYUhyOHFW2AeAqRsyidJXSzN8aHnsfuUpuAiaUho
ggf8Dq9dzRs95uYFbC88VDcgXqh3cPfhJ2UVz6s7dAXz6dCu1XzjSiLzsWNUhB0BRM12OeRfWPyi
Ej05Afmzzi2KfTghm1PdlXO1G9ca+z8fb2Deflnr6VAlVPer1SkckTKtjOPuWwvk+aAUNaA60WRU
s/nOGYjGIroCMjG17ecS0uFbV1H63n48re0dFJQcZckZjgZa/9FACOAX0x6C0pLkxCQbZOa1CnkO
XmDk7mgPQnvhS//7bS80vGu37EsJ62xBGrjpE+18/9YX10Sj2IAg5K9/Xs4rElvxCxn4tyxdMHX7
LpejhEv2+T5QZP7BmxJfCpTMTnj68hSyqyDkmQp9ciHwOtR3juKuUoDLAxYhG75zNZKMz9LtZk4f
74hagaQa0fJXlN9PDJUH7M3GSefK70p3eyIx/T3Q4/ZcCn6Lrsq5Obs4M5YaNvSJcToC0qLU7FnS
EaF4Rd0LE0F/yAX0fIx11xOh8uPTJwPBm10S09G8rjD2JvuHqxkYkjazgkxuRTpk1H5zmp9DA6W0
u9o9Rt5w6wMw11J1tH3uR9Qg+n/Hg6bKLrEOixMRvSjz1QtehClv65iHJIww/XYGbcQ5V8iGk/CQ
wFcqR37RiEQWOQS1tWm66Pr9HoH2j8OICe+MldTAiFG5PN62DvqJuMz+Ep9ZRawznnrKlPUiFEvd
i1Nbyg7jsqTZLum9Uphkts11EJkc41Jay/UA9hvjYr/z3ZaYUPsd0cCCUwpgsnzsp3oc4Cc1SKln
+3GzUo1EfnQaUBhXqk0E1M8MDSkYcD4cY8DrsQ9apzLDoxn5EF++qBHD6EmvBJ44S2QUubXXKj0B
hy0DSG+aAsBsArLt90FPXUQdfszLcMuCEPHwa/rHswZI/7STfEEUQiH7hiJUAt7UdGaPBxmwpoTX
zh7zq9Efl0WORBbng+9rrjLv0YzUzSpT1Zn8gvwNAWojWNUC/jyI9PGmfdL1KR/QBqYBoHKFTVAK
tget1gnvEMo5fj8f37iK0bb+iRAKjCEbRZICARkvTonCqsMy/0omsp8+/G26MzoioZPqFsItrfGp
VOfJerE/lK37Qpg59Te5o3uG90FK7EuJ8/jzjM8SYz+5uzhOtj0MgoLOx0sHVhVFyy7YdPENhkKh
4Odfe0sZdby1ToIxuIRGt0I3BaR6SDO4YuLxvvqRt85h2ffHwxjzB9H5Zv3SpD7LdLOvAZ39M241
O+Ur2C+ArTOvfY7uSc3zVi6hCCTTiTQRoohCN1QzqEdp8ZvxQHRy3aPbTQQvCUQe8YZzRMJINVQZ
MNzPzCMy8QLt8QcGP7qTHNoHqc96cQ3e5iSgn3F3atpW6x3bx7vnER8M7QJidX7lYLlqQmfvS6+0
oH8oGFItshn41K1hs9dfFciSfPO18UkhyPq/1iR3CBEH/mEXlsolU3dE7C+Oy3JXYWqlJ9OVTQ3p
sGS4C3daqDX2+3rDXvVvCpoj4wK82OXn32PWGLX8sO734Vwolixchm2aWuNCPIdHQYPEWuD4kSDg
6sNw69EjQqSz22nidJecLPcNXrQhgD27qt5ZWXzXDBtsZk1kRMZwu11q09gHF48lwtPrLINU7V98
lKtT7vvvSas8sAkt6svivS+Rv50NoomYf903maX6/EUdhSrf5NLogdmS33Rkpe+aMZXCdJC1iieG
3vV5XTktpZ2/dLrFRMSDzPoYI+IhgP8JcS9Xo5uRNt4WCLkEICIVTtR8cX3yClw6P0YNGZuHFSyO
xKf5bPjdrnLUzVhguuz3uA0NLwsyr4MRrg/yJRv2njCQdZgzOU9Qzhtrk/iYz+wUQYXL/Uz6fDVK
sFvgD8VbjkO8n/dK4uSk+Dx5HTZMSQ5DMN5W3pmIyTrnp0yS95bvUxS+R+/KaR+w3hQbNLhq1s+l
NjLSdIGZx7mXwxOi9PwXOsJkYvVaVUq4uxevJAxVByPkjyUGVa7AtG6Fy0AlESFiCs2mdai5TaMb
zhu6Mxdgz1dUGM8YdJe3gpBsBEUqmJP82Vc92FzY11N2D0V1N6+3CPvmnkAzPG4Sk487VBPCDnil
xgGk2ntxMK8r2cAwpjm4gUMxirnatgDo/Q/8uIa3/KZTNVVcAyvJDSknfE8/Hw3RnjteVaGSVZlg
rM9plMmKO9/rEAInNZh0aChWI6ExwsLjlE2SUuKU1f4eAbTerKb/4zzYDseIqzmhbuhoqYb00v3s
byXVRTrku0LrkaonV/5IR5/0sO50aTlCJ7rFYIQ9a9YgfbZ8E0+VPqyJ+Zstbn07gqEeyZKRmBgQ
I9UKwu/pVp6uipfVu/UpwkaO6XdMQhmx5hi0xza2U1Q93ksPEj+XLkQxV1lnWuCEalYiRCJheyRS
CoWft+POMIghcNhrxSH0IKhAOlzaQQjxkh+QRpLj3hVnOHjAejwfOKY1ZajgBk/LRu2coGZg1AnM
lKTMIxisIEEiP5pF2rvbBb1cTPJIM+SMOorKRcukHYAcOstSFOPM8lEK/o42QqLjmUC2Cp+O4UQX
1hUqKzbV2JXx6vHGbOZJUWJCijSGKFZKDZGkxc0igXRHx0ffydveSomdYhJH2SoStxFv8bog6I2E
Brb9W6aZj+lc85jBVYtdr6NVYNPgpsVOLxt+bHJwIjArGR9tGYhIIKhY08gvEWvgBNr6axMPC/A1
3cOwSPD9uFWK0GVGN5jdt37XNUfd9ig+Y0TJkGv5P9kyPWUqml08fHWQa08u0AvrWBdGCgNZCXRC
m5+j3x1/NSKXvSREKQ4MwKQWhzyOFiNFt0PS9a+sVP1Q3S1zNr7wT85qait/DtDD8eLoJMOtZe8M
eJ22C1guecQ4Kz+3caRgTwSGrsDBoMGqqbeSardMylLJXehuIklI41t6JGpOeIJxZZxXyVkeC/oi
JjVMx8KSOBV96LODtlY7Kd9cnJMGcoPtpvBALWz92/3OvxrReJ2knQK8HWy/QtCC3+6F6jYKhNMu
CssgF5l52Z5dAfR0DsBkDrM/9FEU5E8vTYtUVQe7jIVE68A+QeVMsnvfDCImnpuG8PjB0H7OmAkn
2lOPqBBcae7RbA+RX7IdikER1BahoHBoz5/jAuxoxcbFTL/kIYDNMjFBUaa1UFLa3xtHfri2KHAp
OHvCpXFrLLfHlKfnIoSzE1z7918K1kgZ8Fncxs0HPaun9hbmKMMMD5DKRcUkc2JvL2V0pI240R7Q
z2cN+BVOjxu9Igj9190UH41J49Qn/ltRLf4AglAtOwgK2e4Izhr8ooBt2zuYjW0dzhbs0OGzy1AL
c1lnErGgDIp9TjNhouDuxroMrY0RGNeu2umUxrX+6dk9EqZ9wkzRyP/PceB1GlSjMQlyfjRPsmLP
/lsxAgp+LFeW8/t/Yl8s1Ud2F5xw8soItF8nmdfwGlhM9vCwlMSmeo8PZM/+SxCzynmp6PooTWYD
uYvlyQMU9awCF8MWUEYLN5+PaFjAkENxlxLn4vCipjItadsWF/g4+ABVtOkuwVbrcs+Lm0R0+S13
QaHqZcOZ5b7iRl3IWAEkzaj5KtfWEQckBkavBXSulWBJ2UTKqHuJwYwkDjfzR6cCPjVGKQfbhz1M
XFxiyxhaa4asqwj53Tv0HioTgUFlZdb6nB8V5putARmbGMcCLqM43arVcBwvxHDES8fgvSDqYVmB
cMfa1WY4v1YZ4PCODWQDpFVOjrFOSQvHFpFmzek2rr44C0v3nt3p6m9OVk9aWUH+iZd0xnQ5p+kJ
zinQIq9coH/2e6ZHn4HJ50T2oafkmQ873LNl5Ks+PhqPqc29ibGoin3FaQAURU6F53W2Obz3VJOk
9zXTnZ0XnP9T5l+orQSsKLWMs0IMIvASU4ZGoLZJy1bYLu6s52zSxDC9bbTbBhzb5i33nb/323aA
B5bevbLZ6oPVg6hc0Fi5AujA573LkUcz8aWp7FBPwgo9QZkkDN/366D9uP2vjGoHb83xIt1Sd9hq
2pKQIgpFolre0RHgPBwcbtSH9GQ3bap3zxKnHMcg/FhheHe/OaU8s/nGIhyw92t86ysRobQgE2lU
PP1qF5vgelNtuN0WQND6b5t1uY4Il90x2K2J6amNvaHkeJVHz+foaCPyISxn44ukd8rpRSqUF4n4
wle9FsXPrKIiOERYW5uSYZX+h2tMceD1kRkOLWzLlVFqHcD6bwr+hYGicsCawYmIZIqaqxhV24Jp
TGyO/3YHEu263TJe+9DPsMUmG8fjc23YFORAg6y6IBe8XFogWpAMxCKle4uyZyyXBiN2eehD0aLG
lzTzCXg9+cxgMpyRd3XWpQGPhfktChFw/0NSB8Zz7uhawt53ZNxXPS/tGaH0s7HoBgpiu2BswJSJ
BDxLvirdbDnUGhgr9gdbeurHi9YM2FL8Xbn7Wn4+YizpKl76WO2wvelcXW/ay+bDN4uiUnsgJilB
dspxMxQ/vxCeHFvCZZ91mAQd2wR3d+9Ip+Z6kzmYmYEKQaWhMoosi2ALx5/8tX5aHGDBWaEHMRbt
rrZjayl2BY0KW7NYfAVXhbrjvYx6MoTiCm5UX8SAzokjp3ciuZ0ThrczC0Mqx7kc/dIbvoEw5RHL
Ohyr+RlIUu3r5eX2ClHtMYPJj7NOQQfVrAeH3EAbD49czdK7mrX+zt9L9ON0gQCgmh5zxgkV9Al/
3ZEKZhU+iS/1O3ibxYATvMHmGAwNyP6HZGkOreB+mAVy8FpC3/0AJURrMgVEqthF701ax2GPDDLy
YOJvHvhIaT6mu1+BpEb8ZkmERQzMwNkp324wDZL1EqESqPY1zyL1/smXXIKkUwtQovG7DfZTLWcx
lCnYJV7OJDv75gKg1/sknpJfMzRVVuAURhn887ouzo6YQXAgBiSfrexsR96VmwXMgcBAQ4ZlcEqr
MxXeDDa8VpI9e7FsgshIz2HD+5WWzd5hFrMMm8TKkO3yR77SraTSgGrqvjN2ILm4WcR0lWviRpVb
NDw+cY2Gg04HKP1yI6jCRXz3gf9rSkyS5iXllfzm1DD23AAOkcVUc0DmUGYwcx9wd4UXYlQCzLXY
V9pYtSVcH20E1qmMWpKgG5Ak8hGCZVdH8ds/gx1YvEjjR/XbYrNyStXhvUeu7IL0KAbyfRt/sBdk
0m1FDneVmz5xVHAPwe+IcEYPp46oXHwCAFWDhgkXzhIemvBluc6Vu8atn/y8h3TyyZA9NoGXtEqC
v5Gri7CsGdhtcfPEmhbU+g78Q2ETcVw/JgHWOLYmQiIlradiQ07JTuwu0/gK9V4+DhWc3RlFpMQa
55RgYCTJ1f4pqRJG7QyHvFAOJPPrx4xxIUdPa0wYOA50EfaF4hX6hiqR/o1cfONOJB08rv7TcR5i
SUPqWyP6oLzz3wUAFv7oq5sJQEcH86hB37BGLL960HP5Fb6kZ2r6pc9gPG3BKPxGbVBxhkRgSS9A
R2uQbz3+2pw6Tb4FgD6OxrsvSeI6wNaL7k1ZrOyMcw9mc1qPRPgX8dcsxRcM+WFqlsE14C6sbrmD
tZf48zYa2PMmmZGIYC03xLd1DshIohJwDXSv69mS2Mz/4+giC0BNMkALK1WIV0LzApgIjx1+UkUh
1rch5MQ3Ut2zGR6D8FGgKFj50J6L3mUnW95/nUbg0iAq8GgW+5TfKdpjrsibZkuYp1xWExfY+jvj
V+56JumDnsUfK6NsV1LNCyjxt+xa+V4TpXa2YjgBYfQEmpeAt1IKfjAwlC+9HHDzXjsUCnj9O9vJ
DRJ/Bq4mEyRxbtRoJpk0gGUk0snE0rlRpVGE3EQSmvJJvXdHCtP2yPK8v/Z+7593fjV5BFFenVEY
Fa0dDvOSX1HZadio2fqe845g/EFhwXKNFQJ3pSqf8O5KHYDeJlXVu3pCk2WQr6JbfhN9sn1AysrN
+HaVjJs98GyQWreZJNrGEOo/VtzblMsG0B9ELLqAg3woued9r4L8DwWUz2GHbpnkblcJvZ8dmZmg
jpgy9nuTiIbMSQQJsaadVk41G2WnPMf7TAy0SUaKVqTse5g4SuMa6gqJ9+0MZu1ZHQ0c2xrZcgsO
Wlp7BdYN4KBBKNpWUuEyOKx6snPVN5IIhly4pADW/EeNzDj5sITy1WZCa1Wvlev0dIqEJIvEGnfA
gtrTxTEPWxNHe7+Ao6/qFJ8bqF/WPyjpV72dFgOFu5gO8bEnIrEniroiZTN9OduDNxxSPpRF8riL
3dfyWvHO3z0dj3j6wkLJ2d5O9bb7qn0uM+yeppiKeuBRIKuGVIo1EIf2LHNAmxNMikaoRpquB+rX
ThrHtR17xfE2oadIbk+RexgIvAubCgts388REVUJFDzhHNtZjn1KYfMM6HFkSUR9HSd7MG9QuGlU
pEhMA/Kvn6KPXjE+HVKaJXVmJozolYwrTSC3pL5Ps7KYj+KuBy6XxtUhyWz+6krgyxk+WENWYX35
RMBCaOu2yY7g0CAE7TDG0Wra1w6K5Tw9IuRPNNfifG+YUhovXNuEyRiI4HwujPKkwa/TBMdzdGwx
wh/T5KP7fvOoGniY83WRrhcEGp//hXq0txqjK5q+7gTeb4F7byG+1WTMUMV//7phwWFnggVySo0p
r9OO8dwFqColgRhJrWciXacPoW8azCTrGs+1dWKFgT+JcbpigLvijTUNpf6vAV2/T8RXFX2Iwyap
5hGMnmwsqO9ZYz3n+frCJs4zxURWFuv8hm0BLeC/LBNAloLhCApazVQRHMpzru9uT93QRRBsdugD
I/11GX8UBb2SwsKaIX6mQOohRrztiwds4d4wr2brVMFYPeAJ7WhjU5oA6aXI63C+TXqmC8UuPd/c
LdZUA8NuMWlELXgCQgd4yrw0U8Azd7U/WeVyBW3MDmteEWEx8OnUMl8Ik8aCN22O0c2wBvfgxP0l
FcObQgX3Iat73ld3lJLfWGYjPiPhlWzyw6iHfVxcxelrIZGO2L+/KLrhInXqo7GJPAlzrRjogvct
q+laCOzxflDXGQDR5UTlMvBGH0tN/yxgSYpfL1VR7/WSExmKDPyTiZiwhOfrNg13jWkcXLAptneG
9ZP1M/josimmhlZFqlBFEpKCrvuwqbbymNDl5d0e8/PzB/p5foWd5xd4axO2sKBIaKcvPo/JJZkC
zrgm4BkL+F4YCRVEwAqkawRgJnsv6yuESBYzYCbKsyoqjfwm+iq3YM/Rqj2IxbytemRJW+qdFmKT
DV9qrbzrrD8trlgoeQ7KcQE7S4QWR40TYgX2saglPwGwxEh2ocxqtOQc2cFLDdNF2+VyXpSnPpie
UgxZyB0+zcM2/COiqoSeFDVfg0Dz1qAPdx9R8m2JBpTmn/MCWQTBKax736aD4dKZESusHDiZvdTo
W/KMgBMJz4CqM7VTt8tiqxeLfPh1FRW9LL6kLgKSl1Tv0pdbf1CdN0Sq1cdnxGk8JlWnBuuplteJ
HV6+UnuVxcgoteAft5nr+U+oF4aG1LwQ5WiSRXvq7/KYtCYJEIXTjPcIccT9+FCfhsTga9pHs6BS
/FBBKrsrUP2PZfHuzbQ4UKxICEsfWWpWQ/17DweNmR6E9g3nsBGSozkHiJLl+8vSoC5AXCuBilLY
7Lgvi3UH6qK6pkbMqo85FVQllYkl1NeRe9oBqK8+K2aQhZJ2PZhD8aeU8nNhguzVG+6M4eG4OxBt
xPF+dI7uxeth0MgzQ4hO2D2le5n5fdr2uH9/qG4MiEemgyBy4vPzcxGqcgXIHq/bvzqfSi1yW5bU
5HNghT/ltD//PucsEOyHvgLbKy9A9D6grnaUaikRSqG2B9WyFS9rsGKWZroqQ+GJUx3lX7zMihE4
04jK/52yfkmn9SZL2C5syCKI/SnujOKwjQiKgyJOT5OJetlGPXQsbRw5pIPgJK3huObRn++zYfSK
SUBEvpWaiozTLyjg59mgM97VWb1y/70G29QawYpGMg3/XQaNIIfYt5Dm1CtHVWUtaF39UHFsvy9V
EPhjcFzs2sSrMm+cHuGGto25geQwbEgF8Iz3OGpc91louxLNAQ7u+fVdASU3EE4HWkChkTlPn1mQ
SBOTw9YrG/qupJw4n+DAhRjzUJpvPN8T0QEVsOVBq8oWt1HjQ6Qe2iIzoMtlLmGuOT15CncEmb1v
qlzkrlNMG9BWClukxX1CEDObwzb0rMKnLNhgrFvJkSW8sveaSW7SvpfpwTedJK1XrBNP8zlRZ+Je
PbNLsDxe7ozbRP+7N+gYbVxfuk3VhTVDiWetYy15NHUYAJiFOzSrFVAm4IFW5fKpfzfZlvJ0u0Yd
9ufUZx3yut6w4SKK5h0lIs3xMEBp2N3DrxsbnSPiTYX0CTqYhZY071bVCPX3IV1aXQs+J5cogDIL
JnRTqbWaFmFKC6K95wqXk2LjkxtUqtUb4PbeJDZJfzlRV0h+/zQgzOudHgWEvmjnJM5hVAupTxhM
FhoI331++7ghxf018Urd8E+5oa2pSD0UJZffDaiDrZXpCQnp6rt5wDd4npZAT2o6H3LzXUiNtDxh
23pjbNhd0+QbPeoC94pzdNbXwiS9DhBihV2/ht+NlIOQS9Of6NvuLrIejao3WGWQfU1ynE0fu+5j
zYjIod0govl6QM+gtr7fzUGSEZgsI6frrWAafxTmAt+fDIuvvJ3T2ZMn9vg7IM+Y5yPR1oO6Oi+8
7qP5AKBCdvd5Yt7LIBRdPTeeqn1Q5iggoJ0cqpoblX0MXc48FNrxP6tf0J3H82j1WRRzhbIxt/+L
3eUp7oaL99V1VpApU/KXwLAhxQi6qsPW30r31N+QNR01ILSbN4C8jCBUlkVWN2EPPcoFYkGjMjjZ
nUbNKDMkGvBbKNVDuIzyQ7v7hYcn4f/7WGI14JnBt1SaUkO5doMtPgPysQW0be3xuRauedtbjyOg
PQahRVnCusPfehi8/U+lae+mhJVyfsnt7Im27tRIA1bP+MbJ0v05wK3h48KoSAOYC0CnMmgQHk9r
Y4hRW/cQfv4mQQ4mm0IHc3BeFSWpFmPu+vGjlqF7QqF+P9TKpcBs3HyMRzxADlPkRIcax2Hw6z7J
ZtCanXojOPCDIszkR5G7gkRXwSJ1JykQMDYnjDGZJS4/qWiex5Y6d/zoYkCjtfJuHYUHaTSGRyzG
lZc7GFqDkHLnmgL5ok0iMsK+M7pIx5S5e0R7CfSEaR1KqsnqIuqMGbrj0EjRi5RGRgc/iTedkvFl
7IWkQkRmkQyrFkBr/lgtcRrKCBeQXNQ67KLw33av55Ihlfw1k3Sc7fonndjqZPpixYsvtdhvFCOt
sv2uaQeQS+HRQYQMmRxn5qHp2jrlKu6enzyZ5lwNJYWR+REPyyJHyTIY7jUM2ANpEGceTj+HFYLC
jx53Dt0sOMn1b9TtjxKnwRwnx1i3+YF22/gIT8Lm2GZ/dvHRb9tAy6MBs38w7bCz8CwnL5dOWIBJ
O7P6LfnBCEQUXVgrNyxUuKNBUyErGlTQ7ZTKByaw9DFEDmNlz90RQedndwtXTV+EbLcCwtuUn1/6
l9ZTomi21JSq9Cawdm/I7+IvAmbteuNFBg3THyy/zuf8yRApvDq+ACRU2Gf08xr3e2pV5znFvWTn
euK++2XaiJKjU1IHoQRO6Bi/OKhdS4C4MkJiW6a60nGnodT1phgn+pjSbJ35FFeJA7k/Uxhf+cTR
bcWQrvNe/gmFE+81Vej542PYlzumuZivTfoGdtkaaY5KwLReXUMYv4s67SgzJdxc3OcHPF/2S6UD
ZI1P1rPIzX8Io5mCxN2aUySagl/MGtKfkn6DwdLuTNASLHgmPQmTFoKi6k5a9SNdq4FWiChLVq4G
lI7DgAgKDCz/TnYRl2JD5tA+5GMA/Qk92lx1i7MWeVgevB1zEF2KI3sA5LX9nG0yB5+iZD1OQG42
EKhL5zCQ0PrM95YPgQqiXX5eBJonovBBkZ6vLOgZl8uSxfuCuvXK+nGk5WVhngFExe5Pv/aR7cF4
OkJjlVIy65tYpoRiTIIOyJH1VCvvGXiUDlRB17aiUewWuKiDc4t0OXyTZhAmtnlOAarRh5nsel0f
SnAFqoO3ZNM6OkYQ7Qs1Tq+D5nENFVmI2wVOBLtds1aM3zw+oHGVMGBDp4aLmO3NA6e7oGgVVye6
uZRP4rCqGjApdjebFdpnJAanCYqJmTZmPutGS/c7ykAT3vU7o6tf+ZpVdNZzuZdyQyYCfwz4fOC8
OnL5vxWDHEKaf5QOmVH7lU/pAy9conY1MQIVfS6smMLj6D83d41hR2EHIVNRjM3cIHLf89mzRP5R
ITEGBPV11xyDDV8Y/evbNeKA88Eyp5QuvG6xC5k5wila/l7bBcNMgP6vs4azVhm4cvw4WgCXfkqF
ht3e37izCrjWHrgSTWd0ocJgL+Q5sWoerua5eCzvOk45u7UGsOSGjYindrNjc6wFyT5+sXgN/mRi
J5cFUTqMnIGD/NDOQxGnZ9Dl5+RTjc4wDx3hR3kKSl/aLdT1MIqr1B4D8TaeNDgZI/v7IF3Ugv71
LXHF+h+wKCKqJdRvAFGOadDH5BFOELiW/ABbvIOuan/KafxX8+BHLF1SpdxHmyois3aZo4EC8HSU
IgiS901WFV/xJYXqm4LrWsXFnIt6kHdrQ8+8u/ZHC1xJV7Zfzgf3ydFRi0hECX3YR5w4UVJNxBvh
EAcs3YpN48eulDZInP9KbHBV+dR7q5/8icCBQZ63i2n1RcVxG8/b8KedyeK9/Lza4Ip+Amcd8ORv
olB1OOXJP7deRvaAHXvv67mVp0CxaSCE9in3ytrm8RZthjdgGP4H8VZyiawr1qgRmze0Z4DXj4RD
Ybk3+yzRys83lUsr3LgflM2KdC+mm3LvDFEEUC5X41JcdSxrmP3VbBO2mXjFWjwwexVb5f+Cq2x/
mY/B7eSR69bx06eMHy+E184jn2KeAZMyGQzIxu7ZbJjSoE0w+QM6N85VxeRAhZVt9ETY65XyiGTN
dct9TxtELnQEHuLa8sCvDGsF+Z/NNJHfXlCIC9Awcm+cscpm3ZF7llRsQKhzIMY9e4OmqnzyLbTi
TlBnvWj/ozWGYj0IiXMfToKXhynMZavZxnQdgDqyP3oVfBKvYsrz1ItqL/xUDAjJIbCliiV/xeXe
jp8N5KoBOdjicaYmxdlrWum4nYUUU7ynYEsCjV6X3aEKQLfVwey+AKhMoDr8hBE+MjdU+KeuCxSs
bClKiOCXXhaCc+JmEURrLPvE+cB9fUlbSxpxZ3R2vsfndfmBs/Xe9p6yiaA1oUo+uHDgw4jYcxKd
K/LsljWXbnmrT0EAZvIBXwaHnaldhoNW2fL7UrBla8TtWizwabAnR2nZ9jaUNnQZXKZJsma1JzBG
QzNZEe0+Sr2dW3RlaoUz6R3KvDRlI0/4TpFD6LvptvMG9yLK84KVGY4ZTFJ5J9JUrPNcnbh5fV2n
l6R40hVNMwDD+vGFaVvxkrJLfworH+8NDAok0i4mXzHbMrIG0/33JaTJY7stdgdB4ys6sq7Y8C9w
d8pDnxPQdwZMjBVXCoXMsYY5unSLE6quM+U+lTnbr0ir4I/PtiNTGq7GiXmc1gsMu6czu2DB9UBr
JOmZTl9TPZWLzbmHDvJwJ9rv60Jt1u5CpE96axdV0Iga83aEvuaO3P+IcMDQ1WjwvOHlHz0jBWKz
1hZfPfzWM/PcBjAU8eHbDkchdoY2fBhyZr7+WqEBlp0bXJxv5JnLLQXxwtDPAptCijVOij0WYe1L
ZknrVP9LU2imbZESrTtMtbuIchRzZ9kj8wzv+9hjjzTTqsalcfyQkZ1s02OULj6tl9/4qC4oTtVz
ElcGBm5+4rqHShmRRz8CGO+4OYllGT6zUWqJpNvtRveSqhK6r5dfeRcRvpm6KVh6zO1KVqyTVV8t
V7KEbUGorM5G18lTEWKXYcXvrEYtjBINBe0RqP9cam3bLz3k+UcQ/jU5hDS9avGpXMvBr3GzW5sG
Ncg3AZVEv6t1VsCwgn9k9XOp20hFi+v7CTnbx3gsU381ROiaUUsVVCoUCF62ufJlEjEP8Yq4Q1BB
wI5VtIfCHZyR8wj1QUEWRLI7NaLXqwvNnmT5QurUGt7FcFAtR+x7LjdunXYPZlfhFkXptaxKUoDH
WUVztxgoaPwEgYutd3PvD2DOgyv807P7qLgtAnHLqUqcG28DmTR1M6CINrPCSKocOFrZ+SqRPvmX
JGIkvJ6MikpPDmLZdgVdIimSfbOouh118bJJak97MpilXMoa+FpxSixYrPENA7HoQ1K1UwouOUOk
WnX9Ahp799512N1IBbJKIfWl/TPLgyEVZq8GICdISP3mn37uEZqs1HZ85c/6pl+DO0pcy3ok6FEM
gCDIcraet1xuyZEv8VWKZZfqFlGx/F6F9EWkswe7O0MKf2MfXMV/yo1tzN59YjcC6yZcMXpjWWTv
CJACSne+v6+cqoN6zmiPTBmjqB+wIs2Snv4IzS063SKlN78KmQewuY+ANQwq2cd+HgTuqXAWqPYq
RfpIWstZOwg8xPyDuBObc7DHYJc0tKYd7ClANBAovam202BhPEttFgCem2xdlwhiN9xNSXzT2oSn
Cm90pJoJBph87L+RqolPc/xwqlzVA4PPWtOoSBZg8pBhchiDvXJzb2NppTIV3qgjOA8ydXapZjOb
AR1aKUkZZBYh6AOqlew6y0AJ+TL0xdjTaJoUPa5FyIgrvwENmZs/PX6L7TXPmTsesO7NydNjaTQX
2ht94p+V65Na4jgTP44nOF8bXuCMsLcJytvjGZX1ywpzOqkP4LpGOrI3KGRpswroWERkRHYdSv37
kO5LxpUnRsgFZgi5drtqOpsEzVC9CDy1PCeGGEYZbtKAg+EheJkJB+nVCCD503R7/Y7liOeN2TMy
qcLJWcWbOzRw8Ix0iGQhA2tmqxU3cN/kUBwAb2DzPMVd8S94TVvu58Ov54fD+xBo9/Uh7Q8i3eDM
KuvlzPUxLjue9dhW7KoNAI8N8xKe8pBxRACP35iZO5XcHpFt8IMRQf1pUZTlj5CEReOZKPt31etF
+IQaMmEoWVgbv7jHpjgBXQMziqdRZrCtW5x18VMy288ofcDsXu+NhxqDXveIc9T3h3Hph7Vnpr88
xQQyRwMJ2SZ0+m82HHHPoqok3QtooliF13F4dSXXUEM6VbpRr2iOKrFgYTy3sw6ZScmvFDgyYHcH
1jy9AVrw6Ff2/wBjmzXUKUI0ZOD7XWQ2AJAc2qSHRYagLS7zjCSh5XuU90OCjAfvGMbILz+iB9ih
UkoYTIz2Te8yo6Ye15Q598GhsDZfOYxd2fl2+PD7JbFBKGSEQTB+ycmNS4AlXD1P/AwWmmB+Ut76
G7cVFmwrfiAiI1YeUWSO82dTeqfIKqFkV12y+rTe0BVGv7ciTSNgszMMeCBLDhX8OzmwpFaVioOK
/VO/woGdRkFg0DBWoG5eixLieebGpYZiy/acdTynAwC0EyDi5Oo2B7DHsaKjUABkcQMv5UtZPy7V
2B5eiLFg7oeH94jeqQblY7wcTDwndp2xYU7XGJnoI98piIEfLLva8pc2Z4Hw1MCZoNhRTAVmne3F
mrNFWapNYQD6E4WHjIoGGeW2YRgxMlmNLWntJbYqJitrjDoHvoanRyZslo9FHE0Zb1MxRd7THncs
pmzoUzbHBj3IjlofPVLj1YL3bzwzGWZeIx5gy2nyMYpI0v94K/yIuSg2k+/dqp1IRSuLep1krpFV
Wf+wyB0taIJGYGDyDmWlP1CAdHGSxS2qWQE7SF41e7Ki10FDM9rERh5aZLleeVTVo+CicZ6IkCrD
9naEzysA8AG5HdjhPoMZi+aAld8t5Bo9s0b8KAu6KfkOJRwkvjxsnE8nnksTuRzPByhNw11zZY91
cApVDsi/nOn7j5/94wvAZN2E91Sm12miyg8B+tSOjQzLzky30YMlIbyG3pjnK+lsfNfi01l+Ib0A
rqc/xLAR+XlnWVDqyDWMAaT1qokULItXsltqewVEQOKbnPf8jg6zR5P+ESmNFk51Z7OHQgXaptcc
89+Q779RH/RJHDcHrH87q37BgMYcMyz3PozVW0qvkmHuXfnyZ7oO5R8T8eMW0YDcRCbO2ox3/1sh
KSbzQc9GTYTjKaYx79n/QqbTRFXbQ+pMasnx/TH5X1V8Euon9/OwmWYwkfHGXXsfKcyZnYVjvc1X
hs4EnJwIWVcHNs3HyXVef/2/TFoJ7zKNS9Ph7BKOyAx/k+yD7Hm9n5iAml0SQAS3KrRo4RJ4SjkL
q4ZdKXaDr2rGcvlA3cyYJAgOop6iKZ9LIyvxzJkB3Jzwm+vtgIBGGNynzKHG6eF9oFXdDIe1akuQ
QYClTx8l/dtdEvXAzsnTM+w9tKIyMVn6GFx13H30NM86RA5Up8DCyBPoRPtXcmW+TjuM6BnP/JmW
AZEOyznKvL6G8B3Vc41UFIB00z9+Ll9tTzASjT1ejcSsRUhjzlANP/kmN8UxfQUXqxUSO/tVp5Mo
o3irrnIJyHBSiEVoBQDF6YgRkO9oV1Cy+J/7ogtiPJ7Wa1lfKR0bTNvo0IXGiXBz/VGf62KofthH
16ACkanN4nEzGvmsDl+pMn+UzdFrn7DPImkvJ568IAeSdULNX+lTF5d59UNtx0+Woqysxe0rLH48
qyc9T2d7sMCJQFewiYBO4jvXUqnLmKF3RBOP8s0nSLaNmehi3ROKXhXps4sgTluaXl+HjvrBGwYM
I8PzL9sVeADZ75nKViLTU90F6D8ChIMdlOeSwJFtRF7cdeODj/s196tUk0l98JVlf+VqorXn8ork
numVOUH0XkxH1QErHtkhMUN2hkOg0laoo8qV6RVu7IfOgILLQ5VMo8cgRmDZimB1MXTZY+I/bw1Z
7ar1LE72yzMX8FLVdApntm8gMA7SOeexxc9u+y9Ry77R6LkI6QHZfYSpEfOJc+DuQELcskOb1ZTU
bSCXG4dC6Awp0KNchjBptpDvoqyfi19MCF4W1aNKQLgHZeVrCClyhBfuuTOLosLbDeXrKaeIWHZp
y2w9y+C2j3mK4NNATxCXj6Q/88s66OmGfbfqZ1Nyc2oHXJ3a/OLQcxPjnWMUovLcHdx7CFM8msn7
8x3SZRyHsBjGSTUALbi3oGjt/V/f0IOcJRwibC9rRc9Nag9BBdoQmtd5bhGqvJmnvoqcj6J9GvQ3
3y8CexWcY0fP6HM5yYFKt/S9CNX2q/BnBXtkJQXZlqF4VHWcEa/OMF2VJp4qq2kLcL4xwVoRAsDS
fVPB9eJ6fzAXz8SWEJelUa57bjAbrHnSHGsjQkkUFZaPMvva+UI7yACcmgsMtl0PFKVLB/hTAuxl
qZNkEFLb+cE/N1JRYLouWrkipHp9OfwnaNdv8OcNmaAqR2+5GeYB49ZYgZYHvy/xhrK03PJp2deh
GHrfnckorDuMhcn0s10jed05OAlbYkL/d3cfckC9SIKxPO2qo803VQQ0XRYYn1+vWH73FajFE+/Q
JJaYP/lL3gbluqFU6m39mvbSarvzLhEizTqcEzL6xmTrT5Jbk7nGH01U5TLlkPvgIBK7/KciW0pq
+0thTBrpydC3dYXoE1snkWbMyMi11em61Ef5kaH/HwnCPr+cMw/RRYsTOUrLQFWw2SUkcnDTscLJ
TYPZZqEp5IKwyFmfikh7rFxbaV8nnCpMnMvMoRYbBCTk0XnxXywRut2OdbSz3GEic1JxqUTlh1A5
C45cWLCIccNXwM8RCF8Qm23Cxkt6ULbELdR55mzAkHgemZDjWFCvDIcXN9pGmRtbQSbF94WS1ld0
dknVMfQRvY3JYFPVlJinAAlB4pWiJpoP3DocbDeIwDN5LyrEfs7AxquyYzJg1ODm2gzJSwP8iBAJ
CDz+jrzV4y7dtakwCGJYugPtkQfDCFC6EuIZU244gOjIHnvMIhR1vBnHi/lDnRX6k5RbcHLtSwRd
z4UAp66R7e6LadQauPxKLGdZ/FnA89mrQ48AIfz48jMPdmWAjFXQGTSzhaLec2RH/T+I+IH6ZVph
eQZQfzOVZS08oK4srqog1ZW508X4nClUrh0DsQp7TtQa/1M4wc03CxxrR16FVmgv6kEI/liTj2J9
8i4a39xjbwnCoD1s+opf8GdBln0eUEPVdjdhLECYurtwUyNDr7WUAdJ8g1JEjk63B75c7lNPo9ql
URJ/ZluahZBYGOir1xLCJAFkNoTLyq5iYhsQj2UnayRlwyGtSy8G34kfhJvQIbYCvPJe6JS60hLd
v0GmJwzRMY452ywNqwIlnD18Z+NC6lUmVcb9bdCDkdUTZoFQHkiyPYfTaxVhWM6w6DNAxquuGw2J
ZqUuli8yHPvk0Fw+32O12KLTTAvZIkvaD9SpICM7Nl9bpp9xIXfvYbG6O3it5MR2Z+MfyOa1Jp9J
U+D9xnfMDyMdzDzCB1wzY+DTc3qN0YoCDUOJv1L7TpX2sCpouC446TmxLs+2/jlJ0MSYbPs0sW4b
7A3r3lzN5Ws7o0jMEdd36SaFIbGarW6QgugaXTOuwY1WZ6rjXQP2r5jRYIPSQzOCGbGoaHcT2okR
veRifKyvv3auz9UEsNDiapTvFcyGRr5/B9zG/fIiJzP+G+XKIhg9LwAfqlaUzjZg/u7LJzUHCVeT
rvH95g3WBJOJubz4fUdYYM/0DP4Ut0XIW4ir/CLE7CHPFYgsGSZhucwgCpSzYH5JDALrrGcz8ZnC
tSF5xQk5F9F4szPRxn3DqWXqkb8wHLhCyFF7u3Kwizn48/2lucPWcACHejI73QSV3FQXCiwNKoHd
mEbNzQyNt2wjVIJvYpkwsX2XDZmUsmpoIBtg/D8qKIobtRvUAnyTuOQN4SrHtFwMSOleZQK83oI5
E1700CMwN7OTP0qgU0dC+N3Qouxu7CLyGFEkSqQ/HGoYd+/SuW04Fvy2P40RJH9d9srJMFMoPGUQ
GUbJQQ6wO3kiT4UeZqpP5RhMhp0Bk7SAzpfxCXAp9FHpS0zbtThoW6TxmoGHAuL4wjDhO5k9nVMh
pcKAm9lUJLY3ECBLNcqkIBnYy5bUKoRKpsODg1TXQdF8Qs56E1AnadP/BqR0H9Z4LWRp16A9oxfm
J+7uUcNUtVnzAAWgNNyiY+0GJPKZqYw/jpT+Z6YDPBSfMTeAkmWLbx0ZGrFIqUP6T7/BMF0ZjDyU
Yigwbe1Sa5exnvaHKCKofrUw9eQ7477bXfGBdt216KlqJ9uzSTPN8PxDjZN17ggfrMNuinnhjcsQ
jfjYmuw2/exWZg0bR2sss2OIPLA4y6owOhTQ+AQxvyj5l3O1HNjqIrBNsvjhKqInf2RvOy0mP/4o
LbwNMdlU+rR7SAATlnwKmIBRDs6SJnJfWI5yIJnFqrP20nKz2h3acI+pDG6Ax5LU0atRbIkI78P6
Awhj+7Bo7+b1WY7pjSOW6dnOmZ6cXqboJUeGPsTEkJ1Y+TargPCFyVR5JJdRKkUUUnMtct55bgWj
Jic1vDT4IvdwmWi89hy15PsZ6/idC9VoLdL+f4uA1fniDTbuM+dFsb5SCyYIDaan74BWaRRer9T8
xqIQIHCXTh6wKAkH0jadRZ56uFvNYLyDSK4JBuIePkTtC32BRRNzHph3sbgZYoimx174mG6+0/Cp
ydWNqO6YwZz9tcgX9+Wr4MY4HTdl4vKb2xwHWapcqno5//kNAggVtcs/YqhD5Kwh+a6bMONk+uql
TJT8FOygV5DolR9MNUY/lMu7o35r3ISE7oi1CWSlEO8XZfTdqIxCShG1H/6iMGhEQ96zXEX2Nmxa
aeM6sWfdCBoMnMo8C+hoYV2Ax5cfIRnr/JEwbJDouLfpGBBliRqElHoLoAhB/lyg6gW079K8LKeI
UIS9C08bQ9fZ5mxGvie5wMfSDP/hE0ydsoQUkUunAX+Y4EE6Lefgcjtq6H4gnDE9kcc0u2GP1Co6
FAAaF3Fkemt+bk6QJZt7fzfj4b02OiJkPx3E+HihIjNTe57Jw9f8QckoZDEXSIXwDBvfDlv2PoDg
EJlh4u12KmArX9YZVmOYtYg125MGKCA7grstcIwQilklc8jGShvjmw3z7un40jSBe0vy3m/xBySQ
8OA+bDa4lwakQf/TsbtRqpGqRv617VFJCxepwIbyMIDPJHTrgdB2c9FNuRw4OSvQl5EU3z/wG8bK
LXuTzM2X7sBUqnHFDE8rqQCh1C55599xjb/KFde/78wGBwlcfVN/2Y/MgfAqOktvxtOBEkDAG6ra
uTdoj3ecV3NdWPkaeFIUnhjbUvxMngo9nn9aMn5meWJXkkE8x4x4808idrGG63JP4xInMTEItJKZ
Kb7ei5CGkP8PLZQ4lSF9NkFHSZQiY0CoVh+WGNs4959Nh8Xt5Om6xW4wjAdh84dNOCSOy1MU61X1
7gTMOgxd4fC5P3BRv6sDqSpVpeH7DZchGYsI8sNIo6oY0sLf8rkQ/z0L54UIsIxAJgnhNieuBGiZ
tkL55PMXQsSeqC9qNaE209dSct7PP9wUg4b++KcAA2rmT/LosVjRTAF4psQJK9dA46q40Yhi4luo
fbJlqsem4iN9GEk+IXPVeYTKqFtqwXrPQvivpyK01Xqa+WJ1TtEudd6kekXSebI8Zcd3x4qajs+P
rMk+Sc8YZFr1boZMKbednxS/BuoQNiBZkmvb3xtNI/3fxGoK3nAmnX33RtDy4cYK349qzfi61p02
cmVTJYgpDSZQJm9lkxVT+vT8I21BvxcV6tzSe4OAkxfE5LzjPjWE4t4+Mu4rt65/E62MSCQyMgVs
r2MnIj51yyVHhicZ7wJZwKOZUTrZoIqIBkDcyLrAdLiBEpElH5jKBsSb6bC8g6Fw9DhvZbu7quxK
Spj0NjYhJdHPq5g8s87IJBuckjnItSYnj3Oum4wT1WZNa+DpzxBcECJURxnu7zFfjeLH61fdIVhr
515Um2MinUWW0Z6p3TcCHzlqNGjYv9tRzIWlbnzVKZvCJdKq4rT7fgR+kh9vwyMnNfIDZr8gc8ex
liVtsciGzEuMYVkDB7NnGM2JVU7BhTISesrIaxSPeskrvOAMztm8LK1sMjwT+eegY2Nup2Wo0YQU
5bn+DM0zBtvKuXP6j2w4b3Wgk/DxXTih8lZPXTmtUbazojvgRohRQtmo2wodCvpwP2TpFx58Xtym
6Krnic+1KaPKZtHyQ6W8lTr3P0VjlSdB0H05bMlcthWgZAyF36W4QMxqcnEC+doOecdtCO28X/aY
gwGIgbGjRgai6plLIUk3Q0WixSc7Xj+tYfaqpS9aHbLwR1KEeoghIvwMNIlOK2brYTFMTTtHel5q
MWCxjD8+NqV5k/xbk/bX3qNQXdRjml6Gf88nIrB0aV/D+Wwf5nXCf0mF7SSPJmt4wWglL0wqAwI9
wH+2ieGbC1Z86e1c3E//hkdWmQzDGudQLzUa/+x5/9QwygmDo0Irwh4VokCx3ZAnp3jIsteWMz4Z
xWOebgvWsiLLBdTYbXN5s5tMyIxNEOQgTWeHY05eVQRefDOFcqhvrha5s9UtN4Egn4kQ5JdpPpcY
0GjqszuVbbDJ4mX0n372A0dRcQ6L/dC/dMiMWQa67a5pfjCMtJ57KzTj5z+5M+FGIdf0cytFVPgz
NjSge2rb2AINHAq/3Prc5fYTmfRqLqC60+3ur/AWsaWKHhT80F8mzZ1qHYog/mvudIip3iCMU1J/
KgcKNUL074OLyrQAdfuuiiphfFs103cVMdjoa/o5iy+M4C3U+qDxZxBH7WVIwKe5b8BcmxVTGzuI
ym0jk3E8Ko5iSFjC1S9TOLQ9KxTyh0D58p5RLs2XPrg59wAJNlKQKDtWN9GQGxSKPZ8BlA+RzKhi
rTtzQMrt/v8+EuZza3yB5a1IwesvQFpfq3uJCchyuHCI928QsV8gBCSqeQGqkP9xTqZNrpbIb0Q5
KhnhIP5FjQO15B25tXH7alnayi7ykLjUkoFhV60LH4ThIEz8UVgfcsdslWYYUq/DaRJH6feYVp5b
7urkb2qfhAENDs0nXnxGQdUnFgxSwsgFKbpeUhxM8E7hVUoOdQ0pYstVks2/rDLXB2eqOGqy57/y
TD+7I3/aeYu8+89jIUGlRg7idOT7A+BQqyM+gqkQ3B4T+/N+73NhlJ6HxPLglOX2OZUFizRmOiIR
IrvqKO/rAIscLPfXKCiFSObtcnaWDGugc62DMfUBiw83b4VjJeQXnJ+/XKDryc6zvYS8JiHKPzSB
AUUk+Te+YafO/oxBdTiDGSlGNZcm96Nd1z3YxnZTEXw5jIldmBBOMWaaqdSb5e3V4DWMZ2Q9DoIH
N4URoY+Z/IX/6y9+c18+bjveKHBhiOSLcHfyncFg0tfv1Yr138ZeDSuBMfehNt0PHYR86lAbgLYG
pQYdib69qgaoXH6oLzXwCXDIyovEE4+TRIFSJt6sCughd3ybeHTnih80lOCSL025J/xHIOVS7F19
5QUnOrvEljgEXzmDHOzwVDcCA9w0Uk4hsAwFj/O3M3+yOUKc+jcJfX37UqG8Ld7vPBwdWILT9a1B
UqhQsOXNi6pUKpyTBEKK60YeMX5f/+CQi/LODJiJhBO4mKUuNfJW1LHCPbs/48GHVd1MSNYqDm3Y
bp0zG4SxIPfmm/CRJwPNSQOFLMYhWqcPDh5KaWufOrwdazrMyCj5a49uvlbByaVqSImI6GUdW0lE
pHs4l97buPoqvvbtLVCqWzYcp9/kE0dfaRAH7Ymq3o0ZKINn3VwIB8ohPMB8KfdE6WcARFZXL3cC
fjClderK9q38rvJD57Puo2wtX1TdgjqVKGDJv0MvfvWgMWAdKukJgbk4k7vWwiLbFmANbLjt+h9h
J3VxYD/Gl1xl0VVxPaL/0ZkVtAgdxCoz5HUbT5ooRZC22gZpWx8SaJaBXT9u9vF4lb0GKomLKmju
oNLDNfoVy3Rmf3l+tfVfvsHiG91k0RX3SnP8Xs0SFxpjyDtej1AtsUNSzxDIumoECAaHxRjYLq0b
3JBgy3nThSW1XWdzyh1B4RhuK9nPpcTh7ga21iI284k5LI1GbNVVGQXw/4IUJi700XO17N7771Mo
RAXNLRaEAr//8deJXtPazB8pVbuOucpS7TXuGecw3W+YyvEpl+mq4IYt7g0C+AKlqDyuoXEdK9Lf
xxFnORSWqncDbLsNlO6LApVF2gNJbDWrN6lKzdSPrZwpQrM/ZfZCwQ2Yv1j+PBEgkuq3AwiPw6Pn
vF4Vh4A9z6tTB190AUszUiMKNE9q9OuabnZflsNA7mIPRtQRDZs0+PqGgBF9tIwbNld9gjhf5Orn
xKr6ojnhVfC6j23JFzwP6unITiHMrT9Gzrlg/4ms3zzuSWgP6bI2WSN57A9D8ds5k7zrSwyQ8WEt
YWIvQMxLfvpsrvEDS5dcpHtNCtqDSab5X+rdEHXraprS0/CbV6ulKSpOXD5yqghFa78hXp552Pt/
wT0LvIiU273Kkrz1PXAJDc/nWtPhHRLg2EiU/vfYquZmC8ADjHDIb7H/m45t/oZPo8h7v9tDWLDb
uy3EFI5A5LPQ/CVH1onVjx3uDeDStZlVFFOagXc21v60o9tGmJq8rGsMYP7cSi1xrD9zw/ILukZI
L9um0f4Og3Qs79M9OvkPlwT0JM/Yb7j2TZuIfh6XIceU2zqRZC8FM1qbiP3MT3tKWXvQplqKTYpM
3rLvnlVS2xmRmV4z+m3VSvttkL30MlFNxj19g9LoEGMRQ2InYInNkTXyU62gxnxRY+SmU6TQvhHX
4LJbcOrOZ118WbXO1XwVFU34JQxkN6gB6wb35jfI1pLUAoeMGHixObMMTztJ7dJhpfABETQCCG/y
fr7MWBtjpFoeGyNh6up0pGNzDMagogmcX0TQMcYNsQnnFmQeIrx1B7bQimurujFLPdybM27P22Y6
RUuqjo2rIBudlVuFtc3MlakWV67llBgdGIKTlICjxIOzxV76HpRjqfk/jHK7h7U6ltOW/fe20bcU
h6kEx6TG+sAT4oQepmPN7LPzu+SzjHV8tdhdZlmZrQfhTv/pnu9SuY31T2wSW+Pjz6ydv2faqZoA
ypOrsbLHOD7At9GABsEDZyWHPTCz7xtObLdXJsq9urD+x/0dsbNwHUglyLREHgWdeQfj2obRLomE
WMwNolAxIzu/Q2+plEtF1sg3S9TrSbyTzWPt0wPiSVmxB2GGgRLgVU1zM8Ug5zF9tgM4F2DqIbKb
ShaPG7YOeC4hbsqHp2PH6ARhs5N3XWkETIx9VB0vi55uxgBkRbzF9pUFUzWCq3mXJRKQ+DZq3vCS
JNqMgZ8SEgVg7edISmOhl/komVdeUj6eaB8AhUPpCMFP1gaQ29tuXz0TTr+5yAkTO+z1SMvQxgFB
iksFpel77XXF3DtFU+9pMI1/KMHw19vurlGiy2Z42smgU1V6zHSiQ6BuK92NgJqULoy63Y6NhwkZ
imXVm4gK86e4DDpbyPaszqPDwFezOFZszOhcGD6vgiiGFNG0cdLCmSEe+prDA9wMpilUJV1G3mCC
hkpwzCDI2veSncUSHqjwVuyIO/1kJHK8WWPpKygARqo3dGV8NUdefWjcRaQmthzX6zvz0Z/vGD3X
VulhAXpzqT94aN5qxc7qkC4HDpZbNB0RcUeCQ1h0H9NBauQMDQ/zTPH6Si53779TnrOYCvhpIC+C
hTlIz5I0LQ4Hogxx/QUDE674G6FiCThlMUdthPZqOZR/s2+tCSqTqW6DAXZRWLRojzWHJ0g4Tlip
/AqDRmXV16CVH762OF0hi611l0eK0tcu633ulf5GIJfApedS4ygFnGXdu5er+iZdbZQcHlAnK/gQ
oasdVE11AJSYCoPHcEPLnXlKWZ9TJSgyCq9qhseVjROqmYIj+bPw0digqoaLXkD4Ih3bhbeMKiBb
I67HQsUhhhpnhcoTMOtsVFj6xhj/IjJ/5nqWyj2mW/yXAzbJj4rP02PBG4D2X5Fpt/n5qD5+bdDY
uxKPn3eVs6TPbu57O9G3KaunwNVGEFWoAAHkPUnFqpaww6BCQ9fR+NfB9Q2yVaoXE5iMXxvgSYNx
nuPwUKFSxhkckMVoOIoV2dsguvHr0AuShKfVwT99uHI6KQ4BQekMqFQMnZdJPGXZ09ibrsJocAFp
ZGAvG/cFFzrhTcMCJSBqNFlaCzPxNG9Xafk27kQHsmuDD2CFzLz4UtHceP7IQiqTDX9I8HJFK0dN
WTUY46POlPxK3ofLHK1Ckx6aCoGRY32LIsGA2n618TLTo5T10aSdmMTG/2pwe3wb6vne66M5P3ZU
KTuUnKddNmG+3gce+tmwsO/KzcjxJ1s88S4OlCQESTRVcEvFfpENwSLMjnWXpq2joo7ZAvxUzkja
jIXn383Wg29AGxjKRXTQ/UtQT8mUCIAzgsrrhbYVFvL4H2CQjb3dQf6n8XWoreIzagWhrdsC73X1
oqVIz6t1Ugj60KklAQ+ER5XsKF7BcPF4guYQ4XMp4sM03gJoYxBoqPk9sKBGN7T9GO3w5kWDcfcR
M5ZQ0U+1dhBqjII4QfsYeognKqeX4CVl/5DmFSv4ds9yjz6eiWmaSV5ilfpLz9tiNncRvcdfjEw3
rzaiNwOI0LqHWmZMqsMTLQnCD+X1NzY+3BtZ1VnfdsKA2XZyUnfkQhqw2XbGO0bG7cF5SX1tBvDm
8GnjfUniiJ0BEk8fTUff1miXzasXSUjQMHFCQooPQx/PZq5x7RldbHJ5g/RHvL8UJSpEiRXEdHSI
wfQCh8JtBQ15SyqRtQfjcoMyZRsIICStX9i41WV0OREnCPVPPBt4nu/wN7NnrYItoplNsknBTFz/
fc/L++Z50kWlzuz818DOwDG1d2jWUskZKef9ZFVDxe5NmzGLTDqdNQdIeBR3/jYo8ZXPqz9o4qoQ
wgWX7oFOvU2Jspu0Vh9S0OZQrRNbmDQ8PhHGPuOVip9OB/g4KZfbgzh2SYYN4WD9vXFpkytuoDiA
glqNbs2a7GviFSKB7XVfNnAKGH9Fij0NX20ni032xGjUIfC75HSCpFjedReWta1PAe1k8b7aRusr
grj8107I5io4qhkgpPeX6S+W1wq4+wNbQAOifVs3M2yDQLxeOyL4iuKOZGdendqJueGS7M4vQDoM
ESawZOdu2gtnNh0MjBpgrXb8jtaeRnldBejwUf1GUHfOI1+pbXYzmNL5FxK7CZeleCvT3eH/x1gd
vfbZFw8iaHxZDpWoEMOG0s8Yjd+fA8jtFEmZK+V6lU3k54ei3cR3z0LQsWFUBZt1RigiPXX7YlzA
YPq7lIg+hENTG++kSPG2dc86PN4EV/E7Rsj75/R2/81aMW7qC92qNY35DKz6Lgtk21sdRPYmBszk
Z3AeSkSAGIdHVBJU7M9RuWoXFigWeYKte1IV+KKqh3Z2BsmO3UaKNlE9ujFNY03eN2UkMzseg/IG
NERRldJ1tlqfnQfUVIxTnOk/h3UUgMaQ7GgibOZovWhMzGs9vXabFDx9IXq8a8MF7wKSe64IroYS
4UIsKtSjVABEEUQ1WP01kTScBKtUZTZBHB5Z156oahWZ0lAgnTO2WE3OiMcJLD6Q8G4qS5nBkEfS
DL6mOhgL2NkdA1po1ruGcbf4zdXhF1yyrkXWLhl4H74LU4SoQG30B/Rsn6uPeV1PcymTCuuUMsHt
Y+t4kEC08AJugkKzalEiDzNSaT/cblBpaw/8EesQEjYJ2YbLOW79LiOPd90weAYKmFcNj8dBz9mH
xSx71/BVh+5IOGmtshbAtEm/PQw1PFlPjgcv/FBm7rRGQglmJWbDEeso/QkYazKbpjLjgF/3H2P8
Jf7t8RyBoCc6RGxNl282QsLiIbmDxLmRhJXrSIYiTfajKR1EdV2/T+8nK+aXeOvFlO+KexFSebMP
VmhG4bzm4CVNPlvkY3SDaJXLc5g7nFfNNDUBUU3v8RWf3VSvcOrjFCMjvo0GSO8/YMwXKXOGKdrd
l5KeTIEuoUCNOM7ma/vjKKFmwYNP6YZYCXoWaxtvRlkOP/4KRtd5aynDNv5pOnbEL6sv+lTeotOW
5lofWDLOMUZt+y4jlBjf/306+qZfOyvav3CSkmOwPjreO/jYwgrXp2QesvBi0WDxanVnfvGGlG5D
I96FNW67TOCN5zxG7Xr+VI+wfcgwqPe2r0q3sJAsuCJDntETK79xRxd9I9ENSH5HmR/yv44qc/M2
5IlTYpnHDPnTMFcgUNhdKn5EEw0DXBVrEtzYKlYdgyW2Ewp4/W2BshYCauGMhTQiSYlO5LhdilYp
qRKBiGx9W6gByZiTF3+XKNGySZ9cQF1wWp5V/qhKQl946vhmMvUHQhrFc7NZBv+Dip3zHktkrILO
UN+dNYsIy79FgA2INUaIR2biV8QFqtDnvyCr/tIeffYKKQqIGpAgvM7BM7reqH8FIyZKCN6z0i7+
Kpy7FaW/sGILyyOa2rRrF6sw73lmCiI/UuOks8EEKNrZ3PAWDA0JaBWudqqC31EccxKz8/YcrW/D
kK7nBEg4KRNwV9GZSOm7I9oDkLqV7UG0rW1fawWCwCY0wSi3GyW1hHNRSBueutHoDeoRJGFymF6G
r+jQbYF0duBxgb1v4W/HLO63VEubRE4jhiadh5s1clU0Se3lgy4xJsKOGeVqKMZB94SpFxVmOTfZ
uO8ZY+SaSpntGUXcGXboFUpfcxU8nPdlKVnO/MReUgkPCjB6qtx0pMyqqoMKy0S/EwKhbBJ8xopi
SKOYO4zKzDV9F6sYgK94q8xpF5MtZ4oaTpg0BcjIPSFay1IfXQ27D7UULHPvR3o3Mvh3GUvIu0yT
oaAnBaHsB6iEa6sea7KEIhIe5UtsKSG6w8/iThD1AwwK3BpADOnIjqId5owMX7jObm5xj0Ph3iOa
tGF3INx8SCFmCdtTFPXAlsHDn0tbvjoEqUyvmQVkIMyx/E7nyEf7aCqCHYRfIOrGfJEjfZwFY7dq
zxJ61ZRsPEE91SaptJpbb65qAOFB/+Z4WTtBs9bPDcS/ncNjrAs4Y2T2CkOJlhPf1fDvh8ieAnQJ
WWFeZ1bl9GADI1tqW4JentlE3hI4qTk1ncU9yUEKzXROFdsNLs+kOB9dxwAEdS6t0PhpC2Bgtt2u
ZpRAbRUQmM7JGXojVmjjnXlj6y+QUnX8Sfmpc5P2XsEUg2/nYC+F6s+mH3Ihup+JTWw/FAEbf6ug
iPfJGUAiGCzHT3uzJ8HqS3/HeBv+6xAjPGkC0fy4sn6Uxss+f/1BFjldbAFuu19y0lHfbrx1xtfV
h4fAbFKpG+t74zH1QIiVGgOUU4UD+WeMbfeAB9cbTgwJ4o21H5qNSXG0lZLOQ481wOT+d8yt7eQY
JmYkW4wQbiQZEXa9JYNugtiKhsrFdk4kNU30jnlkmhgZ1WJAU5BIOw0F5INC5eSXTq64CeN2cT4X
8hdUaC2CkMuT86DyZKUowJUGkcDJsrFLZCMTl7A1Ux8LlpbuQKEe9nbqRXaW1x0xWpYSNZ+bJMpY
gthLttMRoUAlKSgbRB6wBk+Bi3l23CeFFSKX993pfeZtDceq8ld+RgZqD/+dI00gq/6UED6cBn3G
kiZ1ud8H2NX84y0CeyGIJNYluei1xrfB/yVgN99Z5JKwsXFGDYuKItS01VrYt6dlvBBGaPZ/+7Yu
Tv8s/5lC3Em/dg+4XhabUfhGleAqv+gHqytnqbjUAwZ0kOJ0FM7jDg43T1SHR6IRNewyiBQgUKcS
1dQx00tEQF3mBBpIMcRA5J/3AsSj3wMZu8hdLcdGgt+0Vvem3tTQs4Wr0pDcHVL8QMbPrx15t381
/RhnmB23DWjO3cuSNMtssVJJyh70MfWrg2ud3pnisWRpfxAwIDanq0T5y3RdOsb4CBlZh4L6bbc0
yaXfqLntk8MDvKQ/EpAKuo53a40By/gbbwMoKh+fNaJ8S1Vm0ltGt93mtKqxqB9MUgsFp3HFTShi
bArqDp2xtZWhNnxJy7wRmugSsA4RXwp2O51stGMukCz0cFpWmVg7lXqjdgsc27PQXesRhe+ZedrP
SUkB22joz/VhKzTH6eswsrj3Zru0NkawZQCxW3SCSSaDMmrjlPYvVKOfpuj+UPg+ICgERHwU0WGx
8yJ3j/z8MT/MxbUUlMQuLo7U5/ORa78cp1oYvlxDhJFa4Y1nWmlNxSn7JdD4MBABvi0VQtMwjgIT
Zs68bJ9QlaG4VVH9OBucJvkgy9jxucCJ7fau8vSe+WwCKnKeKOAoef7kUT/+g3vr9wQTRiD6YRKr
7uZyVV+pAB1wFrsDJ3QBGT8rkmiyuSa7TWK8De/2ZT8tr/ahRuL0yH0nUsOhfQzNK2DfR511t2T1
kLMxJmeYI+gbbEYiq4XlHSOkFxys9MtUeONbCbzFSyBg6t+Cx8DlIGpv2XFJX0zwT7BgXEalWeaI
BMbSBq+l4qsCZk5RZcF6qVBqoCNvA7bZpqhF0mlTe9k9wDFCWODR33Ckqf78rTov+0NV5vJd+MR6
XZ1GatMyK2ihe2MXpKs/dlJa00Qv/DL2YU4mrqrYMdSl5Tgs6St3VQwcBX69OlTfH6hlWm4qqAZa
i7jhsETVmWQ66saviMGGIXCm9Wcqxi2Tekv8+lCpVvWozXkEap5oxiIte8VzfWidNHrGoa0NWLVP
J9r9Dda6+Eoqy/65jCX+LtEjAYlVc5W/VMm+XTOEcmzVGQwnTdZjrFRjJ9tjb/6KskfsIDMypxeZ
lbSgEpoaNkZrkdHApo6XJy9EoU36QbHCsL0/tLZntwcFSuTeQ+NU64GBNPdXAwqSFZMeDejHaeM0
Ez8WP7XdZCO+f/ZzVC8ZJG16uEmDP/r+JqKDhJNoGnJEU/AEvlOjW6ZTLxek3eYOBo3PxSE1rgWE
kNz9grOqsSNVYaPt5b/LaZLQUMlw8z99CvcUSilnr6VXvbza259BRf7ulK7pTmO2dWDBPjWqIC+J
OKRp9ndh/CUSUQX3T/zyXPPFPIEprrFA5WWrJcyTmvXeC6vmHaIo89xFeAGuAZ1wldJLhjsH88Xs
LX1fNhH3Nhe/V+SHsZ8raoSKRzfDqQJ5cyWCrrmQ7rEqCChjX2wA4QPfRQnrhVgbbKbPmVk7nmJu
sKhQzLHU05EMFYlNNsWPvqMPeZznFNMpOx0sbpC9ouXFBCAlKcaS6XKuqSjXfL7X4xaRGGcx10rF
dSqYvntlgqgsTzBUBPAxH9siktDvZRM3c+QEvvQMhtpvFT5C5DbX67TqMqOJJOKm4SvxY+fJ/Hhm
Gd1KrVcFDI4bjpOo3QvX1dmSA9smxCsUEn4WG9PHO5DIX56p7WgHqAtBtmwOJJpA/+skcaU1ql06
vwdc3+TER8TQY6d31ogT2dZ/zpUWPSLXONk5IB9kvs8fG4kEsKD0CkVPzdi7GHSK2KfP6b/fbB2R
XEBkWjFD0yiOHc5AkUo0zMRG4qoBBSGTIVtrcSyXc7xuyn5IooyNhasYHxpcVAC6DqffM75t1IFq
8gO2bwgljvHLTpCpIYUSZ/29V2bmUbipH3IVw3YK1MuoR/W+EZS2LGaQkrnn8zhLj/xUXYCSOHIe
s78dqhs4skq1sD8+QkNSHL1CEy7c2fKI05TvXb9T2ipTYUY5M/5iFx3olZ7BXG66BPAUwiCh9T96
3f2w/aaHa1rBLr2Qyc8IeASF46ALrDPUlll8rftGDTsiPgC6YF+/53be1P4o3bTZxqNaFOpMwlgo
81fNrCWi3A929pRLaZl59Rp4WV0xkVpEwFDnftXO8Um1Fl9lxnplxE/Ubwos/ZXfXD92vRnKD1HB
VClOEsZtYVZXEcV8qNjtN3AZxYxqVimr5bjC+/UXcVexxRXwx8Fa4pVeSWriVIbL9Uf0X31dlN0C
uarVempfN7fJsyuC173qiJ83vdnKbHxFxQANfz8IQyfAWzkmjxJgkHj75V6DzlqmfdEGLS4+MSiY
Tx24kLnOAytyUbsvbGFLY187ZF8qfarAnuTmHXq4FM19ESZbSkMpHU0Bfqya1FT8XJXT2Y73mvH2
jIRar8UGqLrC+5vL/QHj8k65kLybDo37Vz9/X8pLrtE26FiH3yUULwOCZuHuJtp8aVSAUI5BoqYB
Loj9q4A6voYezawc/Pyn+UzfIQD0TSrXxoSX0mSivHLHFj6Req8w3jVY3XhZ4WeeliLbx1bcNvul
ksyXYH+MtTocPvsGh6FhYPRQL3EyARpaABhYSIAa7t92RwSRiFsItuJu63qQC/aN1bUGAYkqhQ1Y
4rfb6LMeRC92iwSKdNfsnJK+N9ZTxxyfDA5/ErGqCSzo70dJPa8O4vAtwVmAcFBiiNmYpiKQfAKL
xDICgs2bhr30WjtQVzvOeXNRkEYtURd0CtyFkK1KM4BljfVy/YgZjLRXGgyzcLUwFlMHdkwNTStZ
89B46Q6SXKNez14t2PBUbD3HCl8PJsTHNUW9yWBSXSNIzk9X4NLDtiUwJnFc3zpg2y+LhvdYeEXP
TnfcdtGqdPYYqRwENfiLYU9/d+LdNWfelyJYjo8FbfCM0bh0ILD/Gz4SMLCRZ/yfT9Zy+gK3xU79
2bpM+ZeagRixu5wrkcImQoMRhez9UfanM4gTY2IALj7uRtTrKkio5Tpx92xvBIFcS3rWZLlpv2Ib
IA2fMURAYj77lqjGyWFOhQXlX5Jq4TEdhIHyq9i5dcp52k+HvmV91sxwBN/24MuvbzDvxPKsDx+Z
f2vvikdNSQAYJVLXExzkQc10rmaDGEQpXhSNnGISGDjF9ZOwd6koeh5lLMR3NhwNLkCTsFGDmKUN
mzkOuxBFrScWuScLFpuo046Xb23Hx76HBWJqDEgiCn7/abM+iL8ida9R3iYfwK7NToP0hYrPbBjX
wOwrsHHxO4vL8AKNNbFlSp6On9zZLPZcYBuxz4+o9UR5elQNdzukaVdmzcp8GhFCGQrDekrOOQx8
n8oQqa7J+rn2vto5rp75w5+xbxmaY/PxbwtZ70aE+8iOy6rm0IQVzUcQlJ2NldyvG47Zh8eiUhjg
sUdNJ9Tw1lfzmsrRD5NnAzR79Y90+RvD6V6QLB2slnP1yRQpCCjV2yr1acbthKCislL4msM1W3io
xS6IiZ9Or92tMyuX7YymAzv3J5Huy2YlD4ED0SC0lH+DAvhHpjSO7BixjmhMx+9MPNmnoFKbrXqy
Ya4aVC7Za02TAfhX2rfWQqmI8pzGKvmWvGu7dcsEctuu/CrtIHGovsQj+Jx43i9aLhKpi3Bqkw+I
xlAHenaAQKjcUVaUy00IxHnGtxrqCTCsS25WUmKqa7CB5z+Qde6FAMkImOX8mX8rHLewpi3h1PKf
MXlTRaSLcS+jTVWrv3BQ08F0Qt9hiIgbmqBP/gvt8G6w88Yneg61CBISX8wfcjDlkuIS55tYJe3k
96VtF/xQsTeIAZe/5lV0IUAxZpKJuNLZRGMwd6p23sRUJWVN18BP8i9QkTQjXxG0WWuXbeidMWQ0
zMo4BO3FMR9XgKvfONsKECfOnTcc1YcSPOx8ptqpV742fAwRfA6PnSRYaCDLfyHkXdA2UwbwoOyU
rat43vdFQrCNWaP9nB37e+PJefHm1xLWqS850OIP494ChNXwFN7NlZqyDvZS2gW5HtAuViL4OLeX
pICqLRFx0cMjn3jx96/x9gOayoubQDPwQDiA70PysafQg/iLsYoenA9hE92ve9bFRG3gnjeZzUF1
XVjqPoC87+gMO7igBh/hRtk27i8CN4dOmiC1wUDDAGDgPnbLmmmPRkS4LDakChNCZpFUsQQqlAEW
VUjzgAVtiAF3zHw2g2qK2rSuZZ8TVDe9SkWKt/dd4yfUY61B6hPfhRDDYjeDox4Fn8CycRBuIV7e
sMiPD/0kHj7HHmXFWg5d1wauElsrQ0R33/ubbR1AGvY6Y/EBlJvt16WVMNYbPEGX5kOk6QjOL1oX
veqrwCXeUmJ0jk3j7+EFqz2036wdIcPgiavtskXj3LCtf7gTSgrM1G9sVza6R4EXX+v4oTsXLdpZ
W4PznJRWqGUsbnQrVB39/wb3N4l5JTnTUCwYlk4aow+DSrfwXLlfQb8Gfl5kxgkCSR+aTN5TKHf5
vPS72fXDtMfML4gtAzVx19SG3PXTa/QeBuPSpLKXPdm+Y6njIa+XWHj9H8N1z2CB4OARICbJIJjE
/M1OcfXjzTd2fiEB/33p2GVvDCg4dZNzdx/KxSCraAsc0FHCHoKU0MneTAn+YRuJFB0k64Mb+VFY
r3jGIqOplMcQ5dOFBJO2F52q2AP3Vycux4Ui99y/38ggHyDNZTvpjnZlH18l55DBs6hwFcnm3FRq
OO6DvzcQJo286p+ehwKUsggMvJXq2lyDx9/HmdoKhruvhhpRZB0yA0sNWk+Xm/gPLhRDcSPGM0BG
YWgOIWSrZA+ZkpJu/PPewBWfUNUg4SATUDa87iwiFKbxHcVZcMIiixEIadC60gIE+dq1VzvivCSM
LTtkHUCQXhPJYTGhL+VfYfqg3uBaloO2oPY/E5iv0eXPxY9mnBoy+9srPfxoMCcS4kj3mpnR6WaT
V0F014dc2aVlE+SXc5w7GpcBpEbgaXGBKZwtC9k0rNBXh9lU/QiUiJR6wR7fzyHx2AsTo6jIUmED
nQSq8omRPGXf0tOR0CV0UehVxCcXl8VPZ1u26pgotnhYKcNqRb++vWMb/Wthr4ZDAA6X1bscxGRK
us3HXRPt5h0BwqAInFY3fpYdAfdrEJHjAuYJOyr/s3x+rdTEEJkx2wZTujTPNUKjxcvxwHR/5oBE
FeiwYODarclBFZ/YrUW5/WmIVPGDBmgC8BCrUNgCkxQWWAPseVlNQvlm1hpvEqIMKNJNuJsp3jW0
aEaT0Wa1c1c8F0QpAEgAdTMettqrRF6vDvKwmwgAauV6kepFXxEZ8mDhym+558Mygn+KfWTI4164
350WiALPT6bddntqkgbip+R5ETTNyRHM5QNTEkUr8Ef8cqsnDQ8OMn0WrjEE3Icv0RDP+kUBVU8S
nCo7Sbopz09JCVpxadYY+gGA/vno0kv/pMFc+OqBUiFZ2JboTRyFlJXuQ6AjV8qybAg57PU2ZK98
qjSiSuJvLUH2USuc075CNYPbTBbRll4HwCCnE2NQNeP0HQOaRh5DIHvn0nlOVq7iC86GO1bzC5I0
aygRrrxyxabT+reGkmLydZ/KBJ5pIUsRIIccl5SzQlE3RNqYP+UjCFLUNZa3ifHCoL492CLPG6mW
aBbrVjMae7ahH0mVSa2vg+nlhzsiV2n5RwLJNLYaB9wecqbH4BTiytuTNhToSFK/lxTFQPyp+nyJ
sH9dtOg0WBhXmCBcqseX99fSI5CFC0273OPZ2cWZg0TgfornLu/DunH77qXQvCovEbaePf8zj6HP
UwKLymGn4LEdqkaZRyM7ueIvUyKZ0+bQh8whMDUNpX+ZxXP9G8W47MKZc9k0vHxgJJvYiidCexEg
58TfGqKd7jHenqeODL6J2cF8YieVqv5VlOlc8SpaziUJGZpwfhghNG4X7iGHBECZxlxe7kLrbSrn
Ke8pDtdRfnawVINaNVJcHI31JkAZiYARW8a8uh6YlHDzOHPK5MS4yC54RUzwAQeg9kT21bGbvN9I
UvxnBgbE0L7X3cX6fRr595jIdy0gGkkBKsOwJR0D5ygvCATU9yA2vpVvWLxYmlH8lp0joCnJvbuw
iqyq2Dv/GbdiKKUdupNzy5EUnqun8X2ZXMGHR1GIH2rOvU9c4rY6vPcdywnA7N4djAbNFqAD0OIB
1ERvn0QjzvR3k5hvdhD97cR1sbw60mDifnLrSn1WCdwYfHLYcUKzvftKOXG07644bgf8N0X0Myqo
W9lX4hTGSM6aPmzzH/c8MCm0bD7nPwyPo/op0of6f27CU9nTefdXImRV2QSUTxGIGq+YGWGRQhwr
UkuXMpsP/5W/Q2e4NvIzPyRHMojbGKVXBZWOjlXlGTqafdJzEIL82ib6P0fbJGM9UHC0tqcQtfTO
UTJEbPBEIcjs2RZqVZLzOTdBtcJ4gkrR3HMBJ9d5K3GQmElhgFolS9f1DinZ4Sh272XN7RcfugvV
TRZoYSU+nwynrWp/l9Rp/8s4B4sQnD+WbAAhAl4ebB7I6Jxnpmsv51zFHSqQRIG6gBeQSAH98Bdf
0cGkxKiYax3kf0CNrkevscNLoyusBndLUTgqCeiuRUSKoK79umVU1V/v7N+ISg4jdIwPgEflKUuP
L8QIS34LKz6BODe+pvbUThiAkHUuuchbne6IDfhAfXw5eUuDqJqjnEabefHo8kmW0rOVxRdnMjCA
Y1BvWlvJdjpUYQ5fNeF2j9hStbkDNTcJR/80khZDoSUBDoeT4D1YSliVdDCIJwVYfyZpN3mfPR0p
2loxWQAqJwqCT2+C10N1gxuKUgsDDL4iWfSEJ35TmPGyWGNkN52PwoDDE9MqYGwF4PdQqhtS/LEx
lgZ90N7HSbb1cpnr7cR0R9qxpbD1DwlOQCd8e+39cFfxv9T9DPwu8D/SxnKx0TG/b/IND0F2qyK7
tTQa9KGSPB0tucDiw5TwymjPyhWDqIoobBVhnDFMhdDF2NQVWEzt8QkUFLagiZs88dvkGF8Bn0oI
tqiSS1kjRe8JErJYCsHS5vYI+NVJJ8/0RPLlPMzSYepq8lhrIgnUHk56xuJYMS8iYvBf4rywX77k
4+RQVvKnb4a/1gQPAliCChKhkm5d+HEsRwy4BTqgeYUZO6nHKyCyU7mg/gXAJZty1FU4Px0ohIM8
W67KoaTmUxVowWj3LfT2yrSu4wEX4CfmmiZG9HenLdJXa1VbuOuF0M5CWA0cEAXf40qzlt/WYl0p
jIoSyscwuZafno5OMb2aFTlmDJ9QXzoRFNTyCTWvowhvua725D+2UTPtFGr8xAGcVI7tZNnk3jY2
ksT6Ge8qfwVZ+wZpbG0eu6lO2A/WATOPiKzUycC2i3ipzlNfjoSjSTBT5OUPkgoHsG+cTdQ1FcsS
Gu6o6LL4RV3PEeuQo8XD2wwo9ndmsDfGPPFn5nTLFdYkne0GMCNs0NaWs1CvTBHGkiws5JkSzhFW
5Qvp0OmL9ipub8SH6/hnkMC6uG92dFX3Qfo+jz4EVQgeHiQuudohC8VsbLgI3u0yJzNPs6qhsIjo
nwxvMQ8oXzl94F1BEmKP+N873Vv1cPymDTButh+hPrHSKfOc/CXG2FPec52SghN2xyDDwtQMiskg
sBoTlgqe+rpkhSZIZa3nNErSAKgD+b+ZFQhVK3ah7acxsK7PRpTHwDK6LZ1O8qJVnuqzo1n86F1c
QHaCMl5iQOHqWqCsov7gxN8Xn8k1W8sOQdLmoQnldFy7fY4QF4/wi8wssFL8JL5WCEahDW657vqb
BAMRKm3CiOQX1wwOZkG20dl9Oxw3K5ou8sbHl8Nq7KleSUjUPiEv5xO6nYXEIuHlz7BcgU+BaFp6
j6HOdNsO43hJz85hAjvbXJUxcDdtZjtszE6U5/Z844/+EUyQL6WdmgXDB/kcOxGXcE3LvnCyVUSL
AZhCAVch6fD3s0Wfnae/l+EC97VjwJ6e6CPTbbAi16DliyGbJPDG5f+gCO9fEtFMVj2qrKrZz9Jr
Uwp72dSYJ9F6arJH2IK1jlF21Kvdt08cXoBc5dxtqVkSiL797cch66sZYhlWy2EnP5Mc1EQSNwcE
2w/DHI0xIwlOcde7sh3J/DpyeafwROMl/pUWAfu3DprtuQaXldoD9qNbjmIz4/3g9oVOaAyhpqXi
2ElPpLZwL3xCFUOroAALNywuGlsslr46wJiSc4iB7uY6e0UwtEgtE7e0zhzhqAs4u9rvTlcUK+KO
TXYCPwmvS5IIBroFwCObnxlj5aLfNVrfJROJHlXla1LuvRzbsxEnPn5REHwY2i0e9i6f6gHXa9Cz
1FI0E1mhrpKJD0jOx8c5YTNoi4mReQJOXpgbG4TcgNGaCRzAoG2RiDLo5ZOs8er2LHzojKzxUamQ
ejSJ/8j0qHSR/ZUk+A3WE/4M7gwL1u33tqpM/1BaSE+Iz3/RlhKWbIOHpsbRgxjwcsti73gYVjcN
h/fw3g+o8hziCb/cIiTY9x+qDoayg5X2QBLXadatwLyl8ml/X2crAd7Ds5JufWGtuO/gyvbQcs9c
7s6z9WiMlqw4GWOs0BmL8Wz4eqtHKek/rIoNfRjLtRpWXhAk90ATeuoQDgB5LXj9CeHECSiJhiCT
+i3vVT2A9B93qQVdjzbngGIowftAeWiBTjAlWX+hi12JHrv6X1FcCKpCfEIguSOMfEaN49fAVbjw
ibXZhvl75esgGYZe+YZm9cAFcm09/KVfIip6WA8/9rSTAN8Dw1M+C1jNUQyyJdQnadxG7WlBros0
1ITVvdCjzGtJTRbb2nimlRUTP+nLrkemQ+SWnvWkYZIaXmdliwndOwibHdNRcSPGU9JUpNq1py1i
pgfHfS9sitXGTtQsNFrG39n79d4fNvDjUlSd1alOOTxwDASiSahjcSdKrJ0NoDNBqQhsQK9MR8Am
l8hYaztaSUD+habh6EWhEQAutQ2kLlMBdWvwHcolIObW69M4KebPvKwUf1WZ4PLxWK8pJ5pqAYhK
d5j9fnhi/aSz+guMT5O1g8fKerkzqgQah+7fJL/8p1tFzh4LYVlJViMDg2WzmBAs8vsBw+/jQHa5
x5SP9ZZMtHuPXQiuaGNmwhjmtuRZ5Y48AKvu7rSKHuFbFfC4zQw1yY2S3b1vo7uP4McqADicbJ3e
0FkfLcL2Xw86pA/tClgSnivdDcFi8BL4hKBIA/9+ku+H4lNWeJBj+nA10yyINRxoWyDVhka3h2FG
hq9sG3wLhNlX9trR7+2rP9MpvgXvKhwk2+XsTBZlRxkldE8+kSGsQZzW9f9DOEuLSrRgmK6un4im
JEOL0hQYSYBitJGURuxSgSUChcx3ElreRsOD64QK/s1yIM2MwIodEPKMRlKq6e+G+FF7+rRrFbvl
X+gg6a7JTOvyd320DJSH2KWk3R4C1iINh+NOwLwdSHcVMuI4uwxKj4aeHl0sOuzrtxbLemw4sixr
YSLLrHH4JvyuVRa0ZxPYlkvwBm9RM+3vwxKredQtkIKVQhYweh0GHsPc6fbxRcuvVm9UlSEhH9Gl
mRqGLMc1RpIBmBlIbLw6rI4CfxJXiPY6VdTQpGfq7DVuBXjUpvq8tTLBhTT2N8jv0BbaaFf/5LEd
XHA3oGqm8epmVfLRdseaRwNC+QY1NFj4O4VZMODutFVu2P65M78+smdMV6Ibkny0xOlps/izcU1K
8+ZhhkmR/2jZ0p5yIRbkX+TrM57e/7FB8xsLPAsfLZ+WV7c/bJ00vI32rQ9YWATcZxMQAHZhxnte
Egrsuj2Qe5zTCLA4/GlN2FZnWkPzTY/9VhjdYagRxo5KlJ69zi3f6kK/kzXlbOvvZWOWNnF0WZeQ
02Ff+bHeWHvRb6XGECAAn4UMH9huoQUyjGKGmQuLFETuXLErdfsJpAGBrYBRQA+zy2ztDVMwuH6/
uuYKJQ5riRf+2TRiyyTuOWC1qXG75ODQ9W1pJSzENj41Lp1z7TDvgqegl4mWu4BSzM2mMbDJF3Gy
UjKmMuE/xhDIHhCKn9lO1kWQ3kUteHP+5q4gitzSN19ITw3e0Y9hrCKebh21OuXRZXU/PDDS9fnk
bf07h7xg8K4BGZalGQT1mTnc2UaGxQZdOsAjRqnowywiXoR+vRjPXW7oSdgFTuKiquLVk+NZMffD
LUAKv3AqLCSUtR/OqtFLiX5xNuqLpjgFG7L+JY+7Tc5UlLoL+0UwxB8G1jmoJFDd8f0+ihu3sN5h
iFhUE6fPaa2dDBmsBwIBdtlsAtUxMzW1m75HPb3GocqdtoN7yIP0v7U+X/vyXk6YjLiOScFhcqOw
bQN3SXEhivuK+liF46tbpKEYDau2XWWfQgvOsAcWEsXm2jh7PWhweUpaeV67zz/cplfSou07qDCx
sdIwQPdeDsSfoOkiKOCv6hNyKtuPRmtypw0S5jLmC/Nym86uf2uvN7HtF4oFeXBuhFqVQavkGFBk
bkHEBnrd31YRf3D3Dw9UZonmgyinx0mHyCp0+kiGs/lsz4HEjaudh8FUSvyqesPjZTJYxe50iPYY
0K9dlzxFDN8xCpSpCCqVCsO/AJlhAtNMmSOVVwiM22HFnUShExRHiMmBK1vMfGixzWpR49XYAqQz
3po1bz+8/nB9r4DDrmX2jNaPS2rpT60Jh3nguTiBX3sW4hHEEMwPXnrdaDuooLqI15Wlqm7Dz40g
jtKVaPRpFg+AlqTjsAFXy8a0B4Y1LleWra4I3uaeyKz8UX7K5wo/ixiKeR0lD4XNpJH2vaj8hmMM
FeeLpluVEZ2x7iMo34G8Z+Fu5gDtND+ZtrZ91a44PBpXqcohnv9oJcjm5YuY+uaBJ6g03gcnDzyX
eYZjMMRslhuaKezWVu1ny8EowPyo6QYK+Depp1+d6qkDDJk3dcDPUktHTV33tQlEqElNGVsvYQl+
aC7yRmMss0PhSpwYBtMcfvi3csHpju2cAUGxVDoTflzjnmw/7Bjq6MoNKhIJ6mA9if64D8UFJfti
Rb/Mpz2trtFBOeOAJ9dk1+CsRUAGRS+oyb4R91xN/6MGmce9njuZkZsT6eI2rDF7HgwYppDLA3an
ib12WFbzswvh90A9YxFYn12QfLkQcWlZaYmcMKbirA46i5V6eaLtcXtg3SSpmVb1xUGqyX/E63nC
8ITd7Y3UKDsybtRnWqWhgZPYQUwwgIEiAvDxCcJLDxiQa1MD5zuLCKPzOxLkBJHw/1+IoE71vZPa
KEPQRMkMk0mptqZ2CgqUx85yJzeDHxGUbAZ12FlVzDSXSUSw5Y+1W2/62eMhiXisOD9BkBi6iMss
gj04DeNvtLHhqClPeSsCFohO0q+8Wkd2loj5HHyAaEKOg2EntPR+vjrXKbksSS7JbklSLemMXtdu
NEH7pT5zRc2myl0OFP8Oh7A2uxGddxC/QYTQrNVd+c4uNy70VEZkKXJhsVFah7zP82CJ86ULgtBr
uMEh/K0m05SGwTQCpYGDghfdBU3TNOvEw/3J3CXSUnCbiI6X3OQ7jCJ9IKfNqu8FTUS22jLrmqgv
gHz4bItgneM5k/EqcAwMIGMP2AQwmT+64w7oIq2ETw74wBqvvZcyP8ckcn2Wccis2hR6aifmRxFp
0CybCQ3zUAMGv6sqaXmUzjYSex7hJuqH8SKascdWH53ykZqYHxXzyOKAEhfaMoT5nY7mgGDorvBC
fLCp+8dVg4+/Xeg4Udj3bnvNnSShMr2oGjLUKD29y3SnyzV+uVXPgRKJUf7MgV93DVoYAmlauiYo
8k3+FlgeqmsjQe8NH6X68GgPmZMioVURdBgSLshGweVKj8KhkVmSUlVln2fkTLLLuXnkWYeIH2IE
ow5JdCn5AVZ6ziY2EP/cQPMm0nHg7qxQ8KL7OP4M6Fi9SrASoS/5AQmBT+LlmNNm47LmYNZiudp/
LHoEjmE7dR55pC1pNZ1vP3xyo0MPPyXsTmWWmg4WrahCA5CGd5+cjk/hxRKas19c5Va22FdF48md
w+152YVvzVmBRm+cSq2xnaZD+A7wP1wW4RxifdXCYaQ/BIFujfqxypfx+lSzUCtbJ7IWrl4YrDCZ
YfrSF5D2R6w9eEghsSNamFJ4OjkR6dK2NmUPs98dnml4cc0KzLwn80RC3RpGhPZkPdRqNdpZ05d7
KoNVSdfGn6/Cr4FbVMC8llJHf3zh5ZPbspgEv5mF7JZF0Ov0iko8Ny8wVZqKW9n5evEpe6C7s01p
3346syj5LNUTEfWRSBTqw5F4d5zo2AzxIG5DdFXmwrj8ayrZQ/wXi05cjzx9HbfbxquUKbwdZbyq
MPL0OshlmMDsh4bYmTmAcdbVWNTInmKfny7pYnX9Mjq9s0UXIYbsV5bYB65/N/LVM9A1bicN5AiY
WAadIyivVrkBsQbEwuzLPjdOWsimQGWJzO5UqRPnNdaqy0IbSi+RefcLM7SuMUeNVAAvl4Cv2xmv
ZFn3bPXENkigO6fef1BoW+24qvi3O/jfH52JiBrOjXbcB8yNK52Y7eSTFg2tsAZAXPAJ1w5BVuSu
znLWuqnYbx7l3ezvhvKrTADuIKtSgwCjILFNfQO/bGkWy66k8GZQSvEv1em6MrLhYc14Im5AdgkH
2YRpcfMyyLA1p+8oaN3F4GscOA1hxpljg7s3ktLVAUJCSAyWniAlGhaQk83xk4LkcayuIwXsvrFA
+pylZ+fVom1X5NQHkXrEt9iLw+cp5ISC85b15TQpsC5u60UEr1aHe/8dZ291Qbe7B/flVtVQ2LQd
urXjMwjp94zQd92u/kDarM056wACp7cTYb15pBWYKazsbbNa5CzExFBXA8QalWkTqnDv0FOTdSBI
hq82TIBpswkRQbiC7pwMpH//GO44vTyezntgrTXo9UnEwONdGckrg7j6RbO16vn6kHaN8yJoXom3
zmQVTkQQYUn753Vwagay0XXaZIo0l6o5WP8ULmZsI+bLkB2q+qLx4xdoz93x5taoGdvQOimiUY7y
dP2Xm4/WA76F8qSrSLkEUos7eXqDVKEcnW3u530cgxo+fgk1S9XIpCKBLgPiha0Rqb3Nwh9Ql6qJ
2mmInajLYoQTY706AB94rEjdDweYwEISo+9IG8jSZGjhXo7rZ7tr1g9eJMGTOIVi2Y4tZT9HdH8V
eHvS4cAEnn5RXAcNU0MOfG/LHbhNKf2iH7oysn4Z4DGZ7olPENJLjSNI3Reng4gDSrfLJ5E7wrgl
RgFp5RUBBqDDpDduF9qmfqluDApEYOjJVLIYnKgt/XqJFyAqx9eZnzUOZioZlKp1ACS/BzTD7aVW
8oQoL8IkFgWOJmdiBBov6E9hDG2XinIa8XrpTZH8ZXJZtCWZEFTY5AxmEs8fQ1Ktmvf+zbpR19OB
+hdyippoYGRPx/XADNzvdOATTSQDXbPF+zqj5XlKKSak0HpjNuMVSBIqQtC+DmcN2DzO8J56Glz6
kj1n0b3VeytS8V/J2fGR3ol3GndLBxYLQunfunywf6Cm91XDSEA4HWXo4RCGgDXU0KrBAvHKO1T6
rcfzYV0RJW9XwrZa4DMooQ3pWISLtXJcJmrwOOnVVqdF/McMBwdNsNblJtB4euR2iHqttsZh6HKB
GuV8gmlH5w458zDYj5mrnhhxoQt0/892+DLYkolWkAg0naw/Of4v4/5VOd4S4ycc7SBn9WoMDBNY
jE3N71k3uZW+4LT/jEG8MuC93JyoMelynIrK43+l98FREL6D5/htPRkNy86vLX3AyGcffUMwBzqL
zzZIsaoxlfY+WXJ1FpEDidnl3qjVbPYi0V91PWmQS52sRP7kep1B9PcWZ7TNzaBaf0tPyXVqmDtK
zkzaT8iyLdbXq5LTlYfhwlcsFQn5cepwYDXt8HkMq0Hh28oplNP3e0JNJrlyGRfkCcaycFdaeLWc
KUqs4zJQqGtRSjduBzL6nY2AwDydYHoCEtVMBdtUQSo+j/hu3Hodm9J1IciESveXJy8BiqxJNU92
pea+3zvD3WQAcFyTc+LPUa2Hswas+juGrSpCtqxA9siUJd25vfrqd4VzS+ChBDj77xP457I0dpWf
DnbCH2+2u+X1U0RajfB3o/R3Skh2sY/lMMjZxB5FHRK0b3VQrwc4KuiFzLUR37O08Qewih1uTUi6
O2QX4bIabI8JpzyZY8+11yG1zaG3QBt2IFJW25LH7xL0z9saxqBihsgn32q1FhdeXE+bGmEUQD55
Hi1GiCLFyWzVPIZROjguw740e8A1paLbxTbW5RciHd4p5F7v0/JJwB+yHte0F57eeUihN2IkiA8Y
f8OmBLG/b1K5XXH6OXHpYEsLFSapy5/CH4Rtl1PRQFU9ujF09R2FA4hUN8yP3kofJ5lLFkV6UgtI
83QwdapEru4Mv5XNj01rkdpVl18wiiLIUtR+CPu8qt1XMPtRLsfs+8cAyaBZBBrZESXTlF+lm///
Uqd1Ilfn8/fTnnah0JIsj1NuGM4rXW1Drn21qKWR246jZaHnGIm5+XG47VjwlalciiZBgkbyClWV
p/miafOEX5LNxpsLBVFWjjdc7VIIbQckWySCPD2goYiewHLkOn/IqvwRREI8KgyuRQNnutqIF8uf
PmPmAz3/wHmAaCmwUJ61k/z/UnmPrZVSnLvWLL8nL68X1FG6KVNiz+d5hLsesrQb/YNb4eoW7Vky
wbuhYmNfI1Cs6V7ilRa3ftdYrqI8HYld7hC4ada6yCFWlbNMWXbuBymx5AO33Nj7FAL7Us0bod2p
rSf1IezZThByTcSoXmhGZ8TTtdbCu4zSKVFd+hYvXqBY/eANULtCYUaPAxymuCZ597f71FQIGj0K
E5b3UO7tvfF504LQn0cfjQTjABIhNrkl9IJqkUvf1EgHa/+dWxuwNCcTY3S/2sTG/ZoOtOQhJB6f
2XtI4VUPtivAmNjJmtwZ8jXwD28jAhH1KrA2xfmjfPauiQoPzKwDwav9DqFmsem7bRNs+idwrhcW
LUn9fVUAZf7/8QH+DLFc9oG0pTdvxpO6f1GJ3kO0zl3+nc/R/VURD47fKsy4OQQoaDC1GClOUJ7V
Rc/nm0oREuEPDwBnlkAs5sJyf7YORvu7DPYIFQ2wS35D1QvfRtXx68QNjo4yCU64T8i9rRPDC6cH
YY/recdde6HTtuxT1Obb+eiRWjIrvQXerhKHBqmE65XrO3KnsK+PcD2Bz6BW/2KvXNF9s8epnWI4
pCQ93r2LtexYbnbQ2YYMCwbnJL9FrmkshdMLNnC8mh5vudxY7uHOzqIQBQiB5un2kCtDI55gKneR
kpTmr0akBIR2Tbz521LBBC/pz5GRCrzPhLHdeZb2PTTdcCGeHshpObzanF6skLzpndZGxkNp/19R
jX8YFWI71ACfZEqi5rKOoXlhX5K2TLowPzW/G9lCd3Gpte/lUWas/80xFl4ZduQC2XHr8KE2WYxw
nsU4yFy0WDpPKRTiTzqHvjr5G91VChJbhwb1CoXXUYseFrNL6PiF10jmCFQQcJf49K4sbp5aLScu
lf03UlWMGRp1SUYXQyCR0bo4gM5eI1ffp8BXR1MtWoJnttsIuztpglQf9HsMKUnF0+Khz/V0wOga
dQHcbzb9wq1/LfEUF3Wiu6RMU7woF5ghSpLoYr6tz8u2LcLevwR+OphulpjAgGngA5j2haHIs/PS
Hhvc2PtIDLfIxFBzwaGyjqyzaHkFA3/gJBNwlz6Zl0QOUe/TvFz5YIoPde/M6/4MZoLcYEnmLk3N
4llRhfGga+7Nilhw7OmxzHtdvZ8fV/4G5Bh9MxQJn/ij0k3RoHlIbX3IYHt+yUEldxlVXhZiljjA
Iq4gf9Og5HTzA4sQXUgYpLTb+SJ/qkW7Ba2W7068Zcao6FCUiOGTrV+Is2iYAlMysfOWLha6tOhk
LyY8NF9zrzo4G0rCou9IJ0fTj0i+RVHtrXMQGJtwSjml8pSXjcEk450gvWb3/65K94jE8Kd9S1J6
FCbF7SjqnluKwyElezuRFigfTP4kBjXqJBjTE8fzrmh0lPHXRq9tBDMG1543O+mwIc78EB/SR6Er
dGo7MIMIC96wNIz9sb2qEY6VULRMb6FC1zZhR285OtzyIRkw/thiHE2no/b+i04uPhciPQRwO2Ow
YgvQR8xoo9kzB2T6t9VIa4TlTtGlmtzShiyot2iFB4qzj4ZpE18xPH3BsVXH5sndy+S5R2CXYvJH
a1rRWwhY5mPVppX9A4PWe+iSsuVQy1ov7gqUl934He0lJ4fEc17QTCSFdO9zTRkOHVMJ0uUwtA+u
FGn8sqBP7bPT1spDYQqoAJ4iiqFZTVxZckCGsrVhHm3fvGbu8JB1m+uNeD1LVMC58SuRx9SWkPTo
vDC3LeGC/Lfh21bxFrWsd9x8t0nkiPfNylnlPAZcrdiVFpss8/7iNLLmzTj5/0/PNNXuLQqJRV0c
2oSiO3hB+TbCCci+lTqsmDxeW5xevbu/tHGqYF0HG9SyqyVhr4+NWsTOMIwoUrQ0QCDLt6XQBxQx
EYv70ysKtLTWbA3EO6wc9m0vq3T3QYh29fGbZ/HE0exBmm1yONDvO67QqdEtXzc2UX5o7PvH/RoK
YZB8RYGer58RFchmZE+k/FdsvI4WckK1oNNmfAdu2W2CjIl95jXT99fJbn7ac5hWRHV9OV8A4jYv
AbGFZw10kVOMh/EtibyUuBmCyJy9H1++mWY72cqjoXXsDtRqfYPaHVAeKKwdNKncpokegvYG5HhS
6ZJhhc0IfSoTVpoUSTJHl6EMU7bWOgBYgj3ZEUKxNcLI0WUPBQabWOH7d9gwFkzowOD6lZ63mWl4
SCnwNtMAVHgqSDsvnTj7Z4pFljc7F5I7S7anmBtAfs+Y6WbuDraJNClJp+D6uB13nKPVpbQnJPsn
0J/iVDWlb22E9objMPSIr6lcsJps4S8Z8Ld24CcYMMCmE3U/bV5lUFZ3Cp1+J5v8vh+V3TzLmVTk
AkQgXcflvftHI92fbHmB9hqZypx8wh39fqXBk+R9wyT1DVXjH0uY1VF7ZuHkSk4PrV+43Nj5WHiB
j4y0+wSVIWNWMHtarFnTbWXEVSCq00dLc61YCE9gQrtC/zdye/bM4F7urCy/yhE5SfWtTqJDFvY1
8ph9sHh/m2eNpWylDss27L1Hvi2hnOxf50Iy+2kbqYTVKLpnCIFdAlh1cmwZT8ftz/exuL/T1KiG
HS2j9QiYrXfsfPocqVlDVK8hVjWCgCnsMDnHQOlegBdQ1qdbpiXnXNbrdmTt0K/hKrtljl2bcpPa
M/PimbGbSt+2lkpP+J608UMNe3ahiZiBfWJHRu3bJVZ+PTnpMhbFohtMf+Ibl6OOu0hpfs0+GlrU
jBmOJ0aq0P/7rr/vEUHetmfA/5iyw7dwal75l9qj13niykpgccIBL2MRdFwHzcTZ4UZCpICrdewF
sdGG1/a4EAZYZwQcdeNS5v0mKAUTv+3xd6ssi9ODknKshaTczxFKyKQbxxSfcbtgldN1JSFn7FgD
nBAts+4vNb9HvVaPXuXVmb0B0kaJ7CApDipuBy87srPHwiSgmdKcZjrQrPbfMOLogNa1W2Jmnrus
70V2KESsOXyc7EqpPQ7eZcF1+Z/dvf33eww64fLqMkABYF+vq6k2Rnkh8cCdHwHEw7Rg12xd3XFy
uIXdvVSC3rCS44QR0Z70351BEf61aO+M5ZwJTq93GvsGIRaCOvEabvMWvN6V4U7S2Ssh0xDjsAL1
DHqLnC2w7TFWOIrpVR9EoN86hHjxhr0hNQFbAWILfz/1S013VdEpNPUqFYBK+RJpVvIGAgu/NkvL
h4NUEraqxRex3ad9dWHE1NwgBNJkypwva++FLe/MRscN17Z+BqAwpoLWn/Q8Kwe+L71oZxuH0Hak
NY3j+5dGIGg7+RybVmqwoEZRzpFWSO3N2XpzqqMQz7n8+4+1ELuMxfsk1Q5+Uj5LGDkWRrVWIYjL
1qsCv47BmhF4qy/jsQDnugfONHidrmlMDtXcrHHetztE4R5v+pmiOlL4VFOSilhqTF4LuswKe6Kz
i4s7cDKrxbSzEYphbffPs7jqOSiOcTZe6/jydmWWj8BTpSloNL0G5pO8telSXqqPnq2b2SMi8KAF
pfMboTBbL/u6bb9/6o4jye3s2ATZXzrMsjlS61jDqENIlzv/w8D38XrEjlQsakUEMVVktT4bsmXT
DUZBs4wKNQFDe3L92/hMi17atMpX37QZh0Y0kbEnL+38/dXT26G4f35wPCwWDQKTa1YL0GLd+Ud0
7FcNb3HmQEYYyzSGPoo3EAGgk8HE9RyUW6yI3wZLl6I4N/HzxSXMFs2NVrG/Egg6jgq4UXowlyk5
O/0SYTfk8qC9joRdFKL03Br0ODoozlsgTaowBofcbLFd/q0K+qGrqxhBRGOR+DIWsPb5Uz0DSL3c
uecswdZrJOswJ3Zhvwg4yGlXGXLzKznR2b0p91GS9TJsubll1+7ssFbsVyRx8rY4xHszX7rlKS3+
WcKahHg87ZR7dttHcW3bFraQqLSmtsmM1PlhDlezOLPvhzzlp1iLUIaIz04MUAtoY7n4P0T4xX/y
kJFeArkqvBVFK1x2vcltdKCfeYlO7QdWQ681uAkMCeCrjOArHBpEJuDUD86nI6QuD2gbEnWuwzNu
Fu7W9oduS3wvndUtrRXXBtldzYBVNaAfZvunUdiIZbLxxn9YzMChs2X372YSaG5vej376PkTu/0F
vJl2iD8q2wBvgM3OMAOr/gUfiOxqWoi19MMz6q1V2LseKKl0beibasMJot5Z36AzbxZisyRqFUbu
rtZaaLmAPqDBq05uH1ee4n7fAbFAgFPlUi2ebigwQadCfK2GjLZHu5BvzhUfZxKNXmAqph8+8UIW
36k6r4kSXTeGRICspluGckCgmrF/DSyF0QXbcNxva3lZqL7qQuDU4I0fSRcPocy9IGEf3/2e6IZG
Z9FF1/VPJFv/78jk6W0qCqm0516EDwdIsdcJNPA/U1Gb384JZnhPk90qJPqnPQAXa50qbglKgGhW
uuWFKPS9zPpL1qTY0V6M/3i11zUme/VqwQOsDYnby3ouRz7IUlEtdUfVBY3F1HlWqNX8y/PJqQUU
jsyMRV/WwQkwV9JRXsq6UX+fyIe+qVio6Eut7EeU4jQ2WJ8s58sQnqDFWvgxesdycUJh8F9ZX3/N
6LM2CHk1wVeWdDkIYhAwe0yAFS3qu+zV0w2hYTXzWJnHlJjAYkcbFVHDqfAfWuIk1bB6Xe9U1Wwt
3r8yYRjq/bWXwBXzEk8wpaTwPX0V/OqgynnrJEZMPHelqwqD80tReBIALlRq/1ENpiUJOtFAkfTZ
QTLJH3RgotvX0Sz/jwlzhMVIBSxg+9rNQJUoDsIDcBD/+5wEyqterwsi10OlvLb5rsVUVILDYagi
29vEntbEBDUsBSORcmcnO1y3/q9oBA3nE5EWZycO3At1tXNN7qz3h6FfvDnPRZi+lbcN7NY/2Oat
RS0XcnN7Gg+0LgHWONFILHMzQjVD69XfD35hsM5SBbZ/SkyX1vgtgYxXr6JqSSTXIuQRSYCn5G4j
DMnmvoBGyVFBElHSiI7FYIJ0unscaYMl5FTT993lPPnKrOk3/gfLStTS+UP09DACQyqB4EifgxAJ
ex7RkbTiXqr/hapfHBSUT9TzMuxwLpzm+Px4ozUjqDEIXPtKl88aNoyoWKuKl37kv7EXPKNT5C00
XnzI1oSFLKclA3iRct0qxs4hCD3w8+xJ4XQ+6iibNfiC/LNwghIXRFaJPFU/NyFVDLFa6QYpBxJn
5PQ0MnDzCmQzdHT/u8G531bIeUt02ytP/ITIf99RsWgwzE80VXotwenWvVummphxppWA5t5ktITO
Fl4YrV3lSbtlzSKosOl4fUoY3rpqZ/Pxj8Kqz8OmN2Mq23jsO9T3oCGFTbIgmhAuyb+xNwuKhDG6
UUN0V3LvfqtlZhIcRnDYsv6oLv/cylzuWTf/peob54aJuzEpTAVlLvY9xQHcm9rozxvwUAV/USIg
8dcEpxvWSQfA9DHhLIjwuvGxhxmzwETOB0/neaeIUpR1zAgnIJAGca4y01tYu8eiuxCYm9htG01E
LI0fS/2M8Ubgq/rA22zCMIwFCMzfKwaFWdPfyGYgeG5tI4fo7QKwHqVWPk7Im/dpSZMC0Vp/T92A
el9r4mq7O9AM2JPCqWIjSnO7+yoaIKhEcP0Ikwre1q7+UbbPDXcXYGC5luhUUFwGIEGTOS7grwBX
mhyr4K7oEyox+h6Zi1FbE1SJ4eEh/eAdccBU1ZkKUiNEmPU8vUMCOqHHEg/RaQOaT3EvvW0rEAs9
C5G/qP2PN1mdZIrje6nemPHT4UK38QAZHiFELksraiW3GYHfnXquj1dACDjQuxNlHlUuXEjbuA8q
iGA60evZTUbiJJSx+d4aJ34qA3ZkwuvkJEGvMjQKVaEVgdihfj6iVsm6I+Mxre2rbK7OwstA1BXr
1/FHPgStvZfaUcUWc2BcERiApeeyQ2u8DQn9mHwUHCOV8Jv3RCiyA4JUHgU3MZ7foAGtKJfo/+2/
YhsfNJWcVn+BSmmp2v7ahKZzUJxWr4x4ih2lfnf5alblerDjuZV4P92G/+Xlzld7BV4Hy9kyLK5Z
BG66R5Dh65t3/h6p+2EjRNn7NRhdnixBhGPGEGh9dHrRU1NzBH3IDXRW8QUZDxTA50IpIBsbZKjR
SVTl+XUfDz0ScxNh6Ud+vpHtBGD88EgWS+5X/FFerDysGomvl+z+wKgkSLqJH+oQtO69mm3xvX2P
HD8ZjpDOzFHQS7d7T+JH/8qbEI6v18a2Wd0Jms7XfzZq1DOOLPGLjxJbFSjhzDuCNEp/vqVYEi1K
0ogpTIPB3iDad5QFod5e+mi6m6Jo6m+9Q5u2BbFYAt6ejjAkk8dylxBgW6FgnEnQSE0K2xrRCO1h
T1XWnjQqZUXXJZoieH7JGObcLJkeoWO/cmaW5cJiBZy3Alee0dwFkC74avtCM54oxuUaByT8+UZ9
e8a+tIECJm+d1YuQu4wMaJXOUElhirPqu63SC1sRCJ+0w62vVlETuUEVjQpza8TUigI6xGIfOzXP
H2JXmak0NwjOYfFGtfeM12d+VN88+t7JYTkDNrjIMmSSc28dxoQ/k4pceYujDeG9GXaWWM5RwYJS
nlAgDBbm+1eGffxy7iaWNdQ8NkeX1QVD05oIUM7CzQB3O7i/4+LDcWS+H41ly42YGlY6Te6xZF+c
1OvgtmdnAipxMt7CXeuuZ3KYKdt6L6pVEhEkAF3M2xrhp6l8e6+0uY8N+ag7rBki1hCM6tCCM0Xn
qoxHWMNCPrcsCDx2OcxpgYZv834qo57IlzGTY1dDrItX71E+r+RrolY45ZsP2HFtOQVMmxzJ1qtz
vGhXkx0FFLIPRNyxVooVqPP+6TErSZ4O4ZhfmDNPDYpEeC1ZgW+jqBJr9ozi0qVQVhQflgcMFvki
fzOP6+U8SwmQRLNfaGnE6n3xsJsGAFOXzm5BE3KKenV7N6M9PPe4Cw9mEIwVEBZE7iX8FEkvEojF
5W8D3iVRW8fljCgJOyfpOvSqv59g9rlrJ8UNo5khqOTq81SpdwsPJwEbKwPWflxwzfPP35zhqjvQ
+4yaRhVfip0WpBvbu0tEkF9xCB7qWwIv2zx6qEdf+ZaDflhp3WZIfc2XwtFMCetYXBpBovDx5v46
qZgnJFjGI9mc0mtIRYvRexBHSmfS4Lp4FDiM7GfzqsdimtZUcMM4Nmt60O8U8IxSlr6fpcZhVbeX
1B1e9m5uzHni6x0PF/H0tbW+I7nAlvI3TYZN7ohsJfcl0f43GH/ezyrNZz21qyo+y+KH22uaNBGz
s7U8erM4BWnWtgvd8vqEMie1x6fayKLXz00ZEcgKVRzjvz7P4kIj59ERnQrQQUe7GehRTzFJVJW2
oRkyeVcw9n9qTgDo7uSkv9nHppk62t7Iv3e7VRhmJWG8Pz6r3G2VIJF68jvvM0qIJYLzttc/iLts
s5GmbPJhQiYbH2lmYgb0+pWAB7nRcjZ95Qx2PAN8aShWeQ+fXqDUdNE6EKnoarrVnqV1jtvDTjlS
t13rWq3ygha0nUs7GwUMWmiLZmSHQRhQSw3Bl/nUZAUfc0POjjenByzRyDxQgdGlms0jarDqx5dF
FaYarJBo3UlkN9+W2N3YL6gq8N+gD0MbisoJqm1rqY4jHEv1e8ZvdsUusI0Fb2xaXFIoXUFUt90z
V6/eIufjp9iUKQa6wQh5DtU6AAVfXknRo5+6TIUONRcItE0hfWoupiseGsZ31njurmgPRm6e0YkT
Ol9qzMiQqo4ZvES0KcV0+tlYlAQYliwsnBTAkEmR8VfuLuY8QB/Z48CPagpsIG2+srtcoiMMCYlp
TyqbEGrvrmaK/C5ZAb8HIzhRj8oB+hdDtmQieNeBaXenBZK8k00JgJuOC6xTNUvgD1rCTghT12Us
+VO62/tIjZYU//8AO9/rI4IYYPhn44ey+LslrVxTYWWmxllI5Ft/CpWPF8VrofXe9VaQTnRUXgwi
H6P77zNsuq/lSQ36tAR5COZK1tslHxMonw1zdiPgFSGnMb8yiRTeoXKZTvgNMubIvOcZTv4teaqQ
28nA9AEZJE7nJneV+YD3ELpm5Bw3PY6WlC82LixVdNtaUCCy5stvG/L3diBE1xHBP7fiDXrl2EXq
DiqJUqrNAIIa4XhyIju2uMsp26z0jANNK9ETwJb2hiSzcKsuK/EPDC2UjYdQsxWqRvVIOAH2d12u
GBKAgP9YPoFo5yDKaH1ybiB9Q/W5FPgRM8f8j2Uobw4bH2yBA4sJy7TACpvv1YdsQnZC5X6PGCV3
wXOcknzNo9LnW4WuqZpLsstiujWrzdU5OqmL2a9XVFKsHYJMbeXdYsZKIbHeu/zDSsUGkvvxzWcF
swaOvd+c2HO8UgAVLZVDg4GYWuQWug4APIDXE0u6j2QdPqAnmXoqPCd+YLvnVtNERt5xb43RWaz7
/lhF9JZik97MrkpixucAGB7O5+9VdKOkxU+Dk5/hfLHjsF36KEQR+X6XFiPKeZaXPYff9htvlYn0
kUEdR1UqN56Dn7O/HZNUqg6GiEe5i9TefvK4OAHjgeal1UyjLn0B9NYj3Lw2xLI6C1U7Hwhw0Ygk
0Wz3XLq1nPiNAPxZJOPN9e+IPwSxjZvbdYfGordlZfMw6+dQ3BbdIRjHx/YW/XMzNJgKPPCAr6pZ
xww3QbUDlAiHH5STA+M9YwKPIKjYI2VfM5DUe+VAbj6QRq92pRv1Ty4+mz3qPI0PAWPCUv4hoLLF
Jcn7tfIgKiW1slq7o3k6/jfe1die7DEPgSvmt/r9A5RwsjJ0ilVVf88fD8AouvcFU7Hy4CZqV9R7
zTI2mI1LaLvtRDdH++QwmdyNBorlY8UeYzBWlCByDusoPfiYQJnkAwSGUms5OH34vEitiuhFDncO
FPoFlPn/vo/zoHsbO1iG6oAKjGGu7hXC9OcOA16CvOMSuDApnDAtXmHcPK+NSRBV7JMDdeMi/SqN
7H+KMJqB22synmbiC0EwMARvV9Q2I7Qx8U0s0r8V6aMQfQGFW+sbTIY4ibUe5+wC5ZBnx5/xHd0E
qkzVoowF6n3mGmF4GNm7Kd6CMjA0Dpfj8R4Wg9zhnoH7t12OUNzmfWkHnq/TmTMz697nSSTdT02m
S0lft4gZK3QZ4/BXN+qOy8eVLJU2e8bD8Fj9khGq2iJIU9wiW4d2cABjrHNTotJWBsSIMC09v+il
5iOeiRaMmQVM3Q6ceqQh/GGsIURKfRlxwp++I11NXbeFpHeqaott6vFptZTTBJkBzQHBDa07PDz9
qh9qFXaQnIO5qUCy1iWDgfrV0sErx85b8ndfFMyYkxficr5wVWi6SbhknoZ0HDJcN4swlw9r+BJv
Wsi5KgiTYPEwwlAX4lRoxkDc4mJ3zSa2uU2M2a47JtRI/XSlX+QG1jnsDrV5AN1rYcZ8nLsKAkBP
qZfuYg4wPGJ0eObexUhzN8xixH64InIIL8JfsM0TvJliAuycGbUI1vwUW4RICMOJ7k3TDcHskGSM
wf1bOF+vlDnZm+Jh+14p1jLnemrZ6QRPnH5/JB7UQPJoPKNUe+UHJyUwDMWjNV6qBfagOWIj2m3D
VXIQ/V8CQrvdHlZKp5lBkZkc7ropRjHec4+aycvyWVY3F6RrdIiYOKWfjZ9TrB3qlAxwZe215Zxd
IJVk6GJPusfWqVW2s0L6X5JoyUHn2zGOUI4KBiJeSNpKLBnzlqy4DDi+U5Se1dO4eHra4dc051sw
0VgBqVZLDB2RlI/6uDLpbX8rtd3+yNEp73l6PpsIi7t0fkmcoK7ux+xDs5LFuli3QaUYRVrxY3qT
K59gfrT/caIdkOOca6NS2H2gvvJgA/AQfe+kHNRe1aiws7W4lBadPLo8oer1zTbk+xuTX9/SrndJ
NKPB5p+Jrs+P2cqguOSZv62mk58QWxo7wSsnrhtpdSVuEn+UsRWjuhLxlpqzakP9oYigOuE8o+8x
WCGAQ1WzNrVILm4MY9bOEqlCPe4Xl8JR1SiWbLAR5/MEaWxtV3rQmalnl/bFM9L1nTkLGuB5cUja
5r5rajS55tKWzjcUwhUpDNUPtDPQE8ScTiYG7Afieb3TZkoxpRtnBEADa0Zo7PtCMJL94t3L9IJ3
fFsBFRUiksB6+926+Bmds1SwMNN/5wgo0TPotJSqg8WSi+ohithXPgMDMxQ0DdaZU3r/E3kkOr8S
qGTPfhmopGRpE1DurhancT+xyDRnGQlk5IoteddTfLHiMXjRnaAq9yiOosE6zlRPDJbszCap/4T7
gufmWz0u78DXkXU7xPZWwvGxAoQhkuIZweT2IuLt0Fj1d5/KU9ZWkl1EM+4QA9vbZ/Sgf9u52YL+
DDCMJmFacHxn7HfSZbyXE3PXw5SVyr7en/C8O9ga2yD6R7fjwSXIenGFxvJBb44KmMc7P+W2VOMd
hbuLaxaMHxD/FB5Sp4/ewn9DKiEbUa3DDgmXXOsDyMflFhkUIC4OzP1Zv8f/Jwo1z9F52UUZzxB1
9tzPk3ZtFBLpFnCxxi8yrwTZ0yDvh1QXEENLwb47F4YG5dAz9wQoUTInlJLT4gAvWlVR5gh3GV35
dVq+12IuKWbwsu+7PtJeXxKU1HsoI9fKuR1Cfvx70frHQj84T01RzMTalcWXPlGuchC+nuT3LAyr
Y0qge1mrdKCDodPUISSqV02FYmnk7c1Aa2K3iRtSaeJfvmuJs3XEYFpAqxTkq8dRVcRHeLu80doD
8MgHn5hNhuJfucMhL3pWkCMAT02+yGeiTlIblzdEkoh1oJDspw5DAD7cMe/D4fVuDS5sX9thG7Ja
ZfeF6lF0YBSOVpsRc8FeQWAPZKSOdHROp13iohWgg1vEn+ERyCYlnkUB9NFI0FxpiJewqpaYHvCL
edgfSh71KLDrL5O7mKBmoDrjGOQGX8VJTmszyVQBicAjGfGVbztFPeu18jsJpNmpTvLNaq4MXNnV
WwgvoU/snpgPfj9kmU/YCExP9m5Gu7XVNb5sRSH/oSKU6EUXyrtD5TpFXwkdwKntsoKPvKmhTCDe
8xUk1HodHL0D3OVyvhutgXr1lvIRz9I3+tvE3b0cYnhZSLX8B6Q+j0CI0sEDeTjUlHAssDAeAehO
FOwlcprOiOeEzHQ2i7ViqY53UMgV7Sdwk/Ljpd3EsUk3u9BhRg8Ly2x0I1w7a7Uqv5QHZU2nSyd2
cEL2o1XI82Eoa9vUqsv8WwHAVn68TUYmiRTQGY7qIZk+7eS9ejoAwEVAPNhqV/d6M5yzXdXJCI64
e6FTMH7R64X6bWoTHmUmn+2/p0v2UNm4aIwe+ozAX5XUGfeXmS9dU9jMRItnOki8ei4yMYHUMDF0
2qQCMhnND1FSr7nvhJVdS6mVhmaPVUeyDasm136ZO0IenSwb01rOx5P3Fx3jbUDrCI7lfTzAAbFM
wOxYLomkLBiUjrhl+huLJzXQzXdzO5flaCRg5t9cRl3bcL9ar37dLDHUFIPiwfWWL1+qnZaB+haZ
SaLc/D7TxZZ69CBPfkW1K45DtyUwjtIwp+D/axhFVToWeAnDi6R7Qf/IYo4Sprek2ij9lVvC67oS
DflfHTrU60GiwHKXnKy2NBxPZ1wUCB5OPoK3TJIhzl/56WnCk0P1T9ZAstndhdlCynbexZgXmlo8
Zb5wZ014Bpn8+5ZQe64quUljzY+mThbcGHXzLfZeAT2bWa6Hh5lMptyiuUb1XSNG995jxuSCkYN8
e/2RMYU2wzqs4VkYlBSRwEED8VyKMrEGGutVa82ZXMXCa9fY49YYf41RPa+eognT/atclpGai8uo
Bc7jCVTYM8jEXcyMfwxohLVnc9GVO0ZXRLDIVou+9Gv1KImBDYam86e5CT4ZP5Z26OmVbr98WGss
DkC0WhmqE8i3yfbQXv9QXWH/ytrg1z9V9IB6/OOalbZ1j5t0F9pK+VG72a0lSTCscpIh6IbeOEMa
17JUmW4Em7GzDNMeHNpHXZ/EqDFzxXb7N1QSbOuZMC+qCmzQrzES51+EFk8d5h/OAntmZLkvUhjC
rJFS/5DLEMl8bgKfoYv0WuByfVr/9QAV19DmvhLDNbDhcfK/dwTjSTmU4Pz6kcrsMVfjHcEM1K1G
5ZUvmmUWQgPoASDNAOWiSkT7HsrzFZp5E19HiqWLqENjy0HegVwWEhv8pCDDf4LJ5KuZH+aaQdGP
hSC3+d/8qk7wu9TUFVfPD+eIqHiUTyTFSwZD/mkykLv72Ygm0wYIcQDGAjCx3u8mFHwflIE8aWiQ
u0DTLbiHkAuDG89TbCp8GqTSFh24gxVYEYkko+zZQVNYN+WC32ozKrBbHNazYdLz7HP6zc44tfK9
ixYyFkyxwPmvPuIL2zx/4n6ni12N97FLjWpb3fuTG5XlvtFsMUG49A8NbD7hPTm9AkhFYow+ffYs
dAVM4x5At2iXttjgwz/c726hz53zVAdUF/aYAUxLwsw/Ie2xiwYdrny3oqAUZwT6I4hcMkb0l0P4
RLZiURBQlL89VynmK59uhiZA3SK8dEebS/aQHibYGPDxVgEZ3b9vf4wwyqhuy7mvobV2AgSWgGzn
Eu/LGQogdqW5NNu0NDO8VknpUQet/81lQ72wo5WN9b0AyWJsKIhNSY3fM1SxPghJmfyyrFlNn6fD
raWNj2jeC+astLZakwwtVCBepFTNMpmiPjscEA7tgZsQ8KoXur8MVPe28YQWIDCsGHku7xRuDOD0
TeKcvtbesyg5aZhUPRAi1B0fPJbvtEApFAxXoNreaPG9VaH7gRnxx5fMTSDgVttZm4ZRmKCFiB8C
Fk3uUsvdmvD560/DO+Kh/7JDCmF+yaMmLMpOpHsiQwUz6/5aIelVH/r6UjENtdLzJzlIW0j6+DuR
00ohgfah2ueMJRg6SRTKpzJZpV+N6HWBZSk0K3wxhg21aCRZf9fpCVs4iATFWjjkhxL5Mn63K+oW
Gp3EAoqIud/yMM2PrWAa3klL6l0vzZ51QGYQMw+FKnN/f6WI2+DzJQ3IyQfm70hxuy/GoV1W/mVB
0bAak9347Pec1yAo3lZyKl7RDIlfZ6xnhW5B7L2/SCPymF6y+3/vHDoOYLugJ6iWzpD228RnsRPo
9yKR7GUO0LWzuO9HsxRXLhM4UAKi3jB0IYeuVynBij7Nc2L8VDmbNSdyFUJa1rycHSm5rHj1r0+5
N4hRWGwdeCN//jHLF4R9koJAkecoVglGDFYVDNYBd/i1VUu5/FLCPW0nZHqx4e4zLi/Jennsd0s5
RC0uaj42uJQfZA9bH/zgGTse0ISZO74bBF36hClVe4JrjmxxtlgzY8neAEFXRyeFi+8+/jd02ACc
pQJWfHgg3wHh92UdH1IAFYA55cKUV5KO9TIwk/eXa5DM2T6he+TPRS+u8SQebYr+QyL6ZE/LKILt
zmg1kF+UM3tGCa25TEUDRQrVNUUvYJa8Y2KCr7IlkzZSXOl1XZf30WCXthEpggaahPeI5tTu+p8T
L1zXmMxjbyXz5FXOBibvIIGOn60gT87VulTJdpegDr9/cclehdx9CnTsSNShfUBwvcsTUiUo6e5I
z5hYCOH44ELhd92LqKLWRgstDBVeJ8GHou5tD8woRwYJ68jOtnIxMiDk3Y/unrpUqkoEl4hEXRE9
KxghkRXh1zDlMFI78obvJT7r0oSadCLvVh8d/3L1CMD6A7tjW+HVLD8rRrKRXiTNbjGOEPr+h6af
nEGgCCsj0vL86IHUF1FlEZBpl07GC6H45SAkkwhlZBeQjrEETfZ3sOxE86Ul4Oe/9c8s/8qlAGe1
/LcM6oiDUyfKqfkVqsqlwT44gFgxltbkOVvH6gXd68M8xtLAQjI5qw4Q0oNyFeGKWZplueqc5hqg
fmkdxBqjE0dQKIWGenBTl8EZJ1erk529AR+3qfl85xtyguicfK/sl2G2EmxuacQ2/LzjMozrEbwB
ypF1936jOqof6+EYr2fiONJT817jaNlO7HzyEGK4BktxLPO3QvsRscZaO8qVZ60Wsdo2Jzh8cZsc
62nU1jiHJD47pz5fH9ghTH6KWcZWmIpiwuOm5GJf2GBhqcJadi65fQvcswdeb6OWMztdlFHAKb0j
X5dVj5MfxxQ8q2w26peJUoTE1AD6R3VIMB/lA3dUH7lstT0OvmpRmGDltKe4c91j+pwuqAe+z2lv
ar4VmdErCyFtgn8R3CSuyPouUgeeF9bUR3Ro2hkXpy8d5ZH2mOrg8vdcGfClSXhhUGcr6V2oXL49
MpcPhYDrQHb6Q8ysKmP7b6e+WYPMI1bwiSWEhFUYiXbzpKp2kLprfzqkNW7CrmaUWxqwMqVx4Co2
iM4KO1Nh/SueI/4Xa1Flv5jpVOgsS9Ne7tMXpdmoViFbaL/v+5fYwPJ5h1klPJPIs91KBNrS+rqw
bZqgexH6gN3kxlEICc+II4/ikW0HlsikB0pfksRLuc26cvxEBtV3ouxf39FgZYTmE2s+HhO6n+7C
JeHSyX9jcGFTnKwdwOZcJJBCryiGGDeBanymITHCnkfVM6/qFWvkny74aIXf8OOq4VZcKe1KPmDR
Wj5f4bgFLcbhYisOBzwMI1TIak9ir6c7H9IK0deFN/fFJYZ5AzKSVmcktEAU5zMlueyINBWsql5A
qfEKiREHrsYnkqVNMnVYxFtLjUHmMDv2UIpsSBCSmGj1XR0986GWDCduxioXPH7KT5wx5GNNzd09
cuFRppYs9MAm1IEzAVqw7Mx0KnALQiuBQBZiW19USsXPtHjMoFpxcjJBICdQ17ahTez59rFWR40V
jAfK0c155ghERo8XYwe03Im3VJ6dw1xkzNeAlxNjSWqZG1tcBUUkL0PbsOHdTNdZn0SrZNICV6gl
yg5adzcG5YxPb9JSHd+P/xcDtV7pnuU0CDYsadooAloaC+j9dbv4yCWklRFnrMUX3s81uzGuneEN
8bNU9OsSLpsQ5hUMufOLv4QFO88rGkXxyQuQ+fJedtIfKYkl+ACfVQgnWNZDtKkXYPm1B742p4nJ
YHGxCWCfjlkNMcB3phgm4OJgFiourDn7L8kCj94NfhXphmO+ugElgPGwItpPJPsPYWYuwWbeCQpM
8GTiBxISW/oXz0tKk1McwcOnuipbjyW/EoB4Z479PHaQR4CJ1eiWMHKFGkzIH1v11UBMCZu1M+Pz
PowU6G3hdzOAuwjSLOcXzkgndx8Qcg78nB37xsO9Gl2cIJwFQJ+oZLQmA/po1jES5x7YX7U5/YUG
qC+RSh+34426x2ZdGdxvi2cPXyhZNkDCeWvrJ9+sRrMtBwDG1AvDQuJIjs3quEgwnQTUp9KrO01/
0z4r3wqCUXgY5WHVKme2xw7p4KjFHrnf7hMAFjVheokdGO1PN1fg44YGukIaeqBicHJPan8f6DkD
OjWfagNtIrZAPkGOz1BND4ekinba2ZTnrruZP7pmj8xd9o/EOaTAvjM30InOuxnJrmfX1H9GplaI
eNQwmpCqclnfetRk2fQMQLxOmRRnf/Vrp0QDXMiFNK4qxvesllyqE5n4Q2RDWUBtpVaoWtM/ZExD
WXMuPm+BDVHeyY2Bx8lHEi2w8G1H36v/wKqM8bxPCLZoJ0vq0wINNDFqgOC4rBSz1+v5OCbZUn1e
mzKADbwLZ/hebtC1yLBIW0ZhqqNEFbCPySPLx0Zt9jbfbyRLY39FVySDL5DA3umFPoUIFFJPQ5K3
s/RQt42krZf0WTstIFPiSCJFoN5ADYpfHlIcRzwJQIOn1tBMskMO4sO+qMLTpmdNIYI4bPTu+su4
aQILIalnFEHd9YBkeXWa7wM0F73GCDqOZaSyc/fXCCHa2qC7Wl/iawPz2IHdjABiAcVJju23zjSx
NvxA6UOAW1ycNC61VNSV9dxLj1RhiJqUHLyomCrzn0wQU/3oTiwV3m7XyUuk8U0h3YUf4K+OlJ/X
cVJmFA8PSKmifUISUMOWAWd/cZDpVlt/b8SVia4p3ZLOC9bBuVwRZMcEQ9i08ry/5rSajiC95c1z
vlGh4jERR5o+fsZGzzhpGXDMFElXYsvwFfx1IZZovD/s01TGQwBlnfr6VWc2oA7gPL9DYq7E4R9H
M8dFTlAX13fqzEkZBCfaKn0J7WpYk4EaHFyYFsmgOPxPm5HhxD4mbWZMD0HWsAZGoNSd9rdbs+53
ZJXptPSmiBG8YbxxExKT2vwo09HlmaHw/a0JdoJR0El9RAUCxNO8bPAG8NFzB3FEOD6bdXB358ri
ytJsBocYv2u04uZLPYxBmEb1B5ph81n7F6dSSn0oFebzi9bW3G6e3kZ65XGELh0CtKZLHNRJYfmi
GaLXYLgKVAKjN4hJIVChfeb356UlbXL+XBl/fhLbh3zOCH1/h3kOqY/GNUcUw+EhkRvxvdj5kB41
aziV2fEN2+UCGhFTJzPujWbJH/5qf6i8KeV1PO9M9sr0S6RXchptgjJxeMDfbniI5uR7an3xJw77
jr9YfzxpBK4x7At/nqDfQDuD9PhVBkEmSdjORASuhksKGXaDCHfQdXquYLxlhx1wIrOgiixVkPiY
WJ+XdggZqQRazb9k9AeqXJbQ9g+N8mlbvrbtheFw4lWkpNoRjPS671u/0HHXdjYf+0+8LgCgpdrJ
qXIwUMHd2WjuUbIOoekzHcYVLutu+vUHeqD+yzPeLtP7IT0Q9+vqSTf7xNBaPAw3OHeT8u7IkhOy
mysnv6y+WYKXHBrWcpC/TAhns3X05i0pXSwhQZCWqRQ6IiJj8Qcd1WM1NnBLdF3aLm50Eeti9Nv/
xzA4RDpgzolDmTGsw/Fv4Ak4DbW133eIjhAhJEBd+VaKg1OkArcuQxE3iJg0OSlrXbYqW6B+lKwh
nMVd1/DtuzYcKPBhAjHTx1H6iQgUkVBbxf35ohbO/eBj8ANPwV4DfnQcbk/5OPm2reIPEccHNm8+
bpqEuT/biVMJ3d4OgM95lzR+bsS2U0Ig48DfywdQoSq73t8t4DFlfQjgA5/oARxFrXNlfaFjqCkC
NhdrORQrcAHeDFu+3M82DmzJk7OGC23poy2aBCyuLQ0IH5AIhsegQ0uX2T5353RZ+uKenKECsc0r
5t45N6b0U2kpmIcBSnMkl6HKJNmfK60daqD/FXhQWLglOTDsfBa6bkUkpq5b5Xunl3kBTsHhp7PG
fd2Bc8ZOTfxUUTyfJ0u8BGKTTCFRW63aaaYJ42kLifOsqp+0UsOVhF+mVjvcLn+1AG+lcAdZBb8F
zZofxGZjGnheEUIxGMoIC7uYRAjWYhXJaH4zdRx8l5g5qxZaSMhiXgMkr2m4s08ERV+IAoUCIaAc
x5xmRyHHLz0GGalmKWtJuQdxSLl1y95HGGySKfEY8J+yUIfz8QXQP8Z2hRE2kPeNYaMj/gZ8Fvhy
ncAV6Z+vLP0+oqOPbQ6clfen+voT9Xbrxc4fCC8LdKPnKAIuZjJa5W5kopYN6xxsI54qojkCY+lo
1HvdnRy5XPIOCGYt+XtvesH/MpsVRgSCDt0Xm07sp4eLc8E4yq64Af1SU+hqVzdJ9yBE0MsWJf1b
IK2CP+QOijSeB/TAgca57bA3uBpiWeqst4gwq+8yM3btjPgwlYafRrz9cj6mF7WvBckFvxj8yYa6
auSByY6jvEx9sWcoPKvXWZnpEgm/FcqlSOSXje1oOrvJQYiHYJdGpqjRG3i6ezis7j565oJQU8fT
laDBCjsyCz7D8IaLZRE2hyL1RQk7Xs5bstvoRZhWf1lyOe+Oobr6a+hg0OSv8o1may8VPf1lL+UC
9n/tKcniazWQdzD2xr1ZrxouGL7xc0n4AqQDEQLeCaGHD4EXHq6jugiV2P46+ZtiPyX360BA2KML
9kZ2TEDSmOqJ0RlrtOD0k8MSgNw7WCoNNNjNAPQbQ7xkRQ1fzD85HCYoSdDlqd06pcCb20zaIPXE
1aK2GKGpkI4m9qXSPZTK7Kb3PuL64Egsmum8v7ZeWzAmy++f3TEyo+Kdo4MIsyDNwfGGhg7otnsc
VTZaYNO9FD05wioUwp0tICJB0OrirAyaunJ5dOSfgiZKhVjnSYZhL0eK89YfjBNtk3/SVixdgCb4
gdhxzWHtx2PuJ6W5vh88duUHutWF/AwReq8N3qooaEIWqhttq2EDWzfEJUMDFv1wSX6p1JNFdEoU
QkolisqB56lIuU0V2MT8akiGDBJJ2wHzjD44DzKxuYpCPCvsfdAxu1Lm9g3VJ7CDn+e0NXU1LLn0
TABdrdYqxZuklZlgVJLpOd2sx4fQKKFC1/Gl6Wvc+jdNSr/+gE2xeQmZWV/BTSyXWY58A24Jt+kR
bMs5Tmo9gJ0YN5VOj6plQrXzcSctMKCnNaxlT7G5AfdPWxcHYllD7c9yi1J2JSrA2HpfpGBQNt19
4Hbpaymu9QBmbKbRDqKdPnXWUIHlxwo6gGRgMiBtV24SiiS4zdDD9XF0zdtqbnRCpX5sDxOS/nIv
4Ty5nKTSt2BbWFQ0tSWsHu250Qu4w0j8leRQkQnbDICgT0ylPyFKwQVyMTSrCaa8SseV7XvGhQSK
LbbAvxj5nvb7jmHjow/QvuMWNX4GSjv/B2oddhgRDXoY3Xe2+zJWvQqNn5FZtAOa/kYs7oi6zJKF
XtpYXLbQn3WF2BGCKMgv23g32gjeDD3ETU4PNCaYE0/TrU+fiuhwMPAFP43aSjKd9xjyc9xP0gbz
ugohsIFgeNmdzHrbxROoRT8PUQhyv31Q+xQio3gJiol2zO/ga2syUhAf3uB9TkT2nLle7bgixOQB
Mi5ZashEc8JLCA1Jm5XGuR3lA+QpOjBuU7mDP8wNd4Pu5ONYQVU90qVPHFFlTwlLCPtPmwyk4rZ3
IY0+jBsurIQdQFWuVnzy6cxm/LWBBKTkFGlL3DqXcwRYi8hSM3+VUdqLPENmQgAN/s1Jh+GYvgm0
AQ28HqjC3PTiNA7LZb1MduqgVOjEiGNqBMRwt+HLlW+0KiPo1VzfM1qIotuvRPcipTWgFDM+fdJe
LtrFmbg/1UQuYOek9usWc0fAdh6apELBci00OzFyEELoy+/O1CtNjLB75cm853XUV/o8ezsWlFf9
PV1UU/FP3abSZSpiW3bNt108wKorZbR50aFJZMEcWz1lmpetKWS0vDnm994oiKX+ibND+t6o/ueE
Sa1gmJMA3Kna+XjHnPblIRbAtgSXxhiR6pa62zCIcwOMVxRgcfYJ/oIRCnXgVaQbrlpvYG9+/XTG
w8l1wtao7Hi35yez5NKbTIFloGR4siob5XWi78e05AJGCqmVPZvCQDFJ7dXlTgYeFkp9hEiB/mlC
u6fKNtJdspSC5VSclVByc9oBZFV35fht2lZR0hsYAqqJvk+iaeWQJs5h6lUrTAb48PPkjs6EAFIz
5rQqE1jOC9KwQsIYn94H//Y7NvvwCcPhEhL0bEXtKekRH9sTrs4XCQcuvWRmUfhtm688ReFHv7dr
v1DYM0OSW/XVG2i5w+5k4vV/J9vJwjTjE6sEBFWRKELdPRQkikP1Tg3LgfT3YbujuWvO8UUxqE4E
w40b4D8H7jbvr8b5ULR6GPFbtOwmYSJSfkrgCeSLjJAJPJwA8qJuUePj/fEM/6fEMDjOe73Q6mUp
X5Uw4xiTKBfJMfxKwxOefs8QIbwQ65hMeVw72lJGVgRSgAv+esK17BbEhZbAe59L+I5iqADChKUm
NU9OiMhpWRqkttLXUgM7UPdiTIM8n/Flu5t2UQtjZVD0pqDM8NkYnU6Hwarum1RvPHDq6koEDzet
CtPbBtA1SXLIlorW0SrlGocTO+DqQyfuKwZa4XUHRFMPoAK3zsI0azmIMbCZzlcMx3plBPHgC7t1
ocElR4ZE/QcwCx1WSTguBpheQHO+jl9Mj6GDn87FXEPN0WBMb8vt7aExxN1bvtmeleNpNAeE/siQ
YT5tkqcMifMemMImXOX+7pAbdGjFNEQaTGPRpiLp5ZCNottQZTKVOMccdxO9aAFcrXG02QN6vdN4
bcM2ZZ57p8Xewho+BZUeL04WmafcIb17Szjssuv/CjSFLFCL3smRbBx3nEMdTgsqFScu6KCDdaQr
UwbOIdyH+piXRZxArdD9rb3Z5yLyMp0Jlm11YYZG2mwLm07FISy+O9xV+1vxQHW54zAKivaubDOM
eBCNoleeNp4D6QKDuCYMkbL6Y1T2V3aA2GsyFQbLyhhlaZLKH50ldMA4ClpI2pDg6z+lwBDOca91
MDE3z+CEGnWzBi0wet5/Y0YRUA8PXL6/vkJuhONr2+0sTWigOdp9VHuMG9KYS5Z1zA59XQ8X/JLr
hrnVvO8tkLtvu33OJngOvomAHbqdMWYf/JUfLWAZL7Ss4+R90hpWXGwNMrgLYuQ1ZmiH1QK85KwZ
+tgxUFqwQvWhxpupBnsRdv+1kNHA/0vyEDFy4H3E8S2/Ev9/MRllGS7EJE04h8Ozgxz4TN2+iyJp
ttJutF7fpfS+XduGD0a+BvOCrC6PojzgOtQtD7F3xD2HQw0XO5+OFRuSSFGpe2BgidM8M8/J00ie
AZZPVQzoOCQhNgQrTtr1dabdyg0qsd+By0lTVHAyS7yxScNlJ0fBLkt0qaJeu6XUlJQHs0QKUC+k
pkmOJEQ1YBQA/pKJ3kCkkf6Z2S0hl+TleOpGkXVzrnz9dKE/9NUZMJru2cggfQ3NGxhWB5JG/HnZ
6IOOF9/aGBM4wRt/nFftBackWQbVGGS5TUbV4mzeWK5Jf2otowcOyU+YmBXM1XvDLc+9qtqESXDH
p4tETeVjVUAFccRT9TpSAt+/yuxkjLztedQJEazNAGPfe+cp7rngZBdjn2+qnyi1K6ls84jWzua3
pbI3jJmwqQtH0kyF58qLbDzZm7H+7Bi5MbiGHWxCLzOWnFiOJDoqDIFCTpd5XIe62cJwA6AX/LUg
T++zwRUnZq7AQ7bK79nfh5QiYtaeR8ol+FjaV0ITCgP6pGaGriuPMlN91vsPaGJJO9s0mZswAbrr
OIqRqD8IBZjffQgrnUAOfnxGUfzvsmnBAL5pi1T/d8F8dQzBVBSNlAlQoSYrAf8ioH8MOEMxbaEP
S0CZOVlcGcPNbGaWnBTZbJP2vLwBQ0usTRS/FF8Q9Uh5+GM6lPWK4EGfUilpTDwz7bNFngiz71ew
w6yhdT9iUwIK2KE2rUfFs7TsK+Pwp6vBPqEL1u0xoxYaxaObLYIwT3QebyTFa0B3X6FF/SKkYnyt
OmhV6adRX7PT4PAJ0Bw9wbHzhzT8eHSGzKatK72u41BFv0DedmKHfwCnYErBrb17sLs5FjGhG6d+
k1IsL3D+pfZRGB0OPFE3+EZsT+uxlBVc5iu1xwFiT7zd74+JFKpg8xQtG0JNcOkiwaimnbwZXvxF
G4/pznhhU54epBiXdQ4+XQ4g6KXv+ksjYUgne6JYQjYD9PHKT56MBLromqHY0oSphmzZIf2wnjQo
0z1cH4flJMKWE7Qap0nP9dZq6kTCJzuJqdrWxopKfzl6fleNHy8RrBkcW/fNE5Cg6Iux5JqBL35X
PQeb3bOKkrj8Uq4obefR2sn8ZT2JKJkkEJ1jaGf1aAhx8AbEIASLT0g+IW8Y8lRLPsy1tum5hFYf
WROHY+LHt5nixmVNNn9CZ4fCfepG6BVwjxkdt1UERS5bHPMBgmx0bMEFu8TPHEc4a0Nk12D+gKz1
J7drVjcp1ZX2cP4NPj1+41XUjOPGMFAclicx6pD6nVKZQwzzXMvc7C/57byv0Aq6CbZetd+UQnns
hItUaEUg8pZU9iAFoulMjkUEplXG4etWk113xgAzgfMmBxTGtcDOXBkHoWos7E3U1R4Jk7suoscd
uolwzVpMstPSHNnX5nj3bv0XCbAZUWPFRRn03fEldhRncMV277Ol/Q/NP5WPlshmsDz0tJZAKzxS
wvkfusFdkfaKYyjTGNV6GBxXeWQDn/24rn5aYsgUEL4mEgs2aRmhMAIH697DVMsuKPogbOWnmc5+
+HeprCCl96in8MsPkO15H4kkcsHCsLVhoQ/E8O/A0iY+jvxUClx7f00nKIU7pPcrDGLq9g3gMskR
2pa5zp/Uwu28hw75TBuwW3d1wiTsEWN/FwZKxVNsqgqCAESjzcPVY/l8N9ujj+JXNeBKyV/gN5GI
6mjQgj7hqA0T2FI2M7C1EU4YZUmbL1dZtSTQ7+yZRx2Eyuu1fXXh3AqVnS9iAe93D80tHkF+FGId
t8hqJ/+fHY6oub7sXkqx31mzF8z1HFrW9dKFzsHkCkLzP+D+fPXm3CHpo88Ykb6ueMGYbn9Spotu
lwSG4muYuY1VhBU/XPSidvQbtUUaDxT/1vHLWaYLjNOXyj+0CNNeU3ugv61TbWqptl4AfCeqgkLD
G0ZS4W47WMfODl7Ia+6N1fJowRhy3mqdEiEhEQDf6bbiiVQ0XwqfFSo5E/0qH+4P/hqniiwuYk5X
9+hZue/O1pBLxSZ/YM/Zpw5POXVjLjRnpS954huL2IZ2UhLPkYFW7H+WMGlTTtzbHNjJQEsru26k
2320V5xppwwdFRqTFvBj2LRNHigcPn+xayY+ydevxyW+x18MQHBWnfccFbzutHHjFWr3DnkfCW7K
rtNtHfjyvuXuCAh2vmz3xIivDenOFCzCerNw/BPQDYKb9GwqsWok0bEKzQNyGVPPU6asRh0cK1rd
s0c+kv7Q9A2hwrxqxVQ3KZwT0OXAE19I95nSQQSMg11q/v03MK1jG/2gW3T44So7eG1U/F49Fexi
+9AYCuDE8XcpK9K4ZClnzLyYWBhJcZ0wwM0EgdDSVUhevxkBDvZsWc68HgzeGDjlLfHmzNcc0MCQ
topO2Q2OVONqr1fnTQ37l3MLKKsqDv2UiqnKswsnLZKAQxCxfHQIf7mRXfkvGKUYZsxionOcwsa4
+n+xGQ6sPROj8Wa0eb9z7swYoYk16ZLYDx/CHvnsh64xXt+kyYe/jxBhcyJgMNA5HprkUGqFCkrz
fb7tog3Ko2HD8H+KzAu/y136Fe8RC0iqbcH3l8LkifuIhCSzQrmBM/iRMmni8n6JY9/twYKtVK//
jW62L9kG5SByW5rkZSiGOjaOAEeTBfW98vDR5ltjI4FxIIb5KmAYqhrn9vWANvOVQmKik0wKmpiX
GBn5bp3QrJFXa3vudg1iG53DwemE5amTbSLCL0BFJTvjAbYKGuz7U//lGNNzzYnC1zPzKXn6mSHn
G4YzV69BKSR/a0kMpHZPJf9nPkRPlf/v4KXVDT5eedi8fd9042yhQVMwysQZiCXwyB2mrSgOi3le
y4O46KiOuQyUJH1XTuXPXO5LDH72bu4iUKpEYoTEbZaZKqCFy1wmDA2rq0d5sTplxbOgM44kBdLB
gYwytGwA1o0ToYVsmCtmdh2JguPMr4brwdEurOioMR4YFDyFjlF5bRnxcxgRPLuGKfSS26lBJb2G
iGaR5TiRarkOrRO9EsAwm3Qaqd4v/NBBFnVOX7CrNUMcMsCq49mz7Tbt80M00yRcSQDLGRDzIZlD
CTWffPp14WsDE2yS2x3nnZMdEHavEXqlAiwyPKJ8nBc3hUvbYs6moQJ1UD19o+kjokxlorzAxiZk
8qdePWNywKcdWo/RU5f63YiQQ5BtHTkA0Hfv2fDUAqQJIJobCWREG5Y++RCH9jHDr7AmNKml4qlF
vB9CV6h8hNPVMhX0aFeLsOc/cPdH9RP9FfBxB3OAq7Dl0JA+r8WxZGTVhxiBMvj36eN+KfxftEW7
vglNe8RiIXIWOAUfWWYr+ixH35ZqQvNliNu/Q2NuHFk2FslzyEpR1Quk16CDpxb0al+6yLimHqc5
Lxkh90qfo/NNQ7us86IUoW+4CYz/jfR+6ErnAXtXQmq2RdI7Q234DzBgqVKv7NAOgP5Dd6hxyQAV
02akk44SOZV53PYP6FGKybC9pYl/YSWj0qIT8pdoDhGf0k8Fj9+w2SNiJIDnc7R/ArQRLlzelaxM
Uj75Uwx7pDX8grd+HAs3hZ1FLlPjxAzLxmTVRntj4rbMknbW6W7atvNp2dbTgkcBGgb/ZrGdfh9b
jyNV+6/6Zg8u1f0yvFO/PO1zHMvAaApSH7X4KwNtQgBsJHp1kWzUjyFzV9PHBEWAyt5smVJA0noc
sEAPdmnBzhrUKwSXtyfodRYam9tctdtwMQPtJzP/I/vpeq0SFQkH8gK0hsl8RJ1vSQDUaC6bVuDp
dsR1lZYHLuccscvvmvs0lh0+C34tOkJ0YuY/Vcyqy1XPL8V8GzZaTvuQMr2KO0nzH4TShhMHrSr8
8QMPn25XRzcNpcvlo9jmuUHiFsVD090L0zFEFz55ZPwEzHMKHKrWAWuLFyjjOj5AXYuu5XeFnv/C
Hp+6eI/I7rZw1zi2UvYo49PKrW9fwcN7CSyWb2Y5jwnF7f/VvVIR6d5BK1iWvDxsks7f339h0pZO
CTyohzMtywpzXxLZSPevgGjpAHSpa9/JCuKbCdYZECCDagqNgeOf0jDuwQ5d0HXfMEtVedL7WThE
8qrQch3wYbbyLmfaA+RFALdPudjhC550fqCFz3TS3obnvMULiO375JzNllJKO4Hp3tNvFD8JJlGy
SBh6iTBVW+M+o+iexCQ2fMywt26UzLniuWtfMuPKHCHA/Kkvtg3oqF0ZwuGFuTFe5Kakq91XhiqX
nKq/GLvhEIpEq7ySLW/oFKb2cX2SGaMyEwdUNf5bA99fofYxm7ijBFl3MhZJL0A+zvS8dBAXwhdN
kZgG1BlF0/JjCTc3mgkT4VsyT1bNcTZRH9ZEvIKPj4yzxv/NsuUEuZV5nrHLymC9d4lxQXkuYcV4
1Fq+9cFQ49G24k8mH7pWOcZpWGPFNWXDjqO2IJ0G6K47xLqzrnMrAplxBY6tPrjxOfWXR334FvW3
q9JGAVZubj4FzE+JcI18+D1LMr214eDRXhWI3/usjVCuRSdOa229rpAs+zcsCWdbbXIrIDecpHLy
9Hu/4rBcQ0pv3HwJE2xe7dn2rmONsDuid5xLEnDk5Hfp7Lz70AuJipFqpybBSwkOMR4EYvkQqS/A
i9jTuBx3wcTaHTpTBcMThsr1+Oizf1p6a2kX4zsez9KKEvmiLIVi/gH60KYocgTrbNA8R8kTrLGX
V9376PXh9c9o0MQ1whErJvpB+uGkgK16VTLa4nTG6A2D0gsLsTk3ti2bBMQ9cqjbhWoIyzI7vxs6
Lf/9ULLSgWxuUoupAV6UuSTM0QMALzszMEFF5uv7ecyDKyLtOsJFXHxU3tReiGhv/in5b+gzBHrc
c+VlnAwnoi+AFgs+RbMJCLzaUKyuf+yy9x0gr878wYQs6h02MvzfMxLOy+08TVA+72bH1tSwcXjP
sZmPnsF1jLao1s5wv9FKCN1bU9aGCNKKczcelffvvgH61sWzH06V9SCJkdYSPCccfu8ylS0ZHBrW
EH7VsXV3LLxz6CMx5Uf/PTqyTmZly0v7Pf8F3uGNYXl4DhTFZvKnfXeYQIQudn/hCAmdoPjbBwcN
oVbliBvHZAebPCUbv+GUKO4eMwGu/JJcvBXeYLR8+W9g59gnZKrYR0UK3scRclGslhvSW3nLNI1W
wC+yg336qkRhGPbExJpguPSWELGZuCHev0U725nDC7m+h0jIcIlRq0DjqrAdEst7GUSDCm19Kz5k
qloIRvJSsJsrmTnCBrodQno9hPathN4wAQFW0ZoOq1B0gw93FYnr9DbSSFj48qXVHHVVTmXb5Lmp
1flYw+0QlqP5AlHH/axzNYeKUa9QZWcAd5qM/K7LPd949a9ybVNgPljKA2ysjtCZg7nWmW5HMoIo
bGUC5TgmG78YtMWO1dNScVd2YYxw3eiN3xaKyNjvUieA5t+uWa7h/06y/j6dLOItnuTrGAtodO9P
YxfX5YgNOT6VE7vQ6RZwrTE8GGo7DeQSx5DZs6zLbKx2pf6/0nECeWhjFwkiBTu6s7Rh7ZpYEarH
BI/a1w0A3Pvz8c78Su6g/fF5DH0c11BbuSP+ib2p2ShsZUx82cNqL7Hro7RgpdvKrfVuQVdhLzzv
ToDhK4JZF6CaZNBvif0MfXQIz8SSv5FK+Y/9ytjcyEe8RHEt/v14Hi6iegpxF7qH39RJ1buD0ZME
9UDzT42wJLNn/3k8glfV5H7Dv6TogzpBmUSjWGdl9KJHWy/NWoVF9SNSKClORTIwbkMFtozKT8zB
9uHhuEmY3wLbW8wLeS1TDoNjxO7TNhOro2CAIkz3lswqeVUCeNQura3XW6uX3jkD4iljQHL8V9VP
YouTHIjZKcY+Ps2M+caIUcIRUqJA7mRlBurJavwcXJ2T9DZwAac+dBNkhphtUtplCJ41Dj4ORBeQ
UeowybUEayAjGuJp7PyjTYXZCDXN2SY55laL2tEOA26M1OgbOewJGlDoJmJ5qh7L4lOBAGIf8w+2
fIgGfe2bYhGyUrsyqx64lnAh+9yRFHYXekOXku3mpL9kBuLp1lIBDWvMjBAvPJy63lJGmZUEIrcx
UFAxp/jSZapnQLlRJJlExggbpRD6MZhgRyc5HbhxuEv650CaU0qmbOgwBGc8+xphpkJpcd6n7KPJ
MvGP71N7sdiw8UflX+94X+gBHzqsvh8z0FAaXjgyySw195zAd/UhKIChB5X8AHGHcyRZL7qKWRg1
VF15Lj3jNRmu6bLPnXB6TEmfUKZlxNapdaAzp8oAXttZ8xVI5ldvAZ6s8LYQzoiVrsdkZCvKkWfo
vWZLFAOlU65PG+G3PH8THVCv5Fg9eikInxIJEdSBC8LEccEXMXTYLo8f9gMEFahps9Abz40bYLCA
FTWtfF+5X3f+4nAw5sO1JiCFJoDlBsBacZhEOlYCz/BhNGvHNf9SSEjRKPRZcr4+VbuGANcR6e5r
9EzlUwXPey7ZQ75l+cJab9PvKW18eVZq2Br4LchAqnNCGrKXSwxOa0GQXj000pSMfK4KVWgb8L3H
E+SToShzUVVa9nRtJwHUSwI/84fBK8hyKxmLnjI92CXakwqtEw+FxJfHoi766oVNeEF9Szte/h7Z
ijwNwGyLCapiEEYthCtDMNU0wjwyKnmpQU3wwJKR2ipA8SHLUxZMaANuVo3797aBoZE2J1hx4XrJ
kcaiwGSKSzrTUq1iNp1dNUQeiamuDX9YVAXVqbKpFk3XIV/Nb+7PXfdOcdZcBsDEO6SNqovFCbb5
j7+wkSH/PNt8Wr4Vx5l97dtZROBtPsmcZRUDn43zuB0Z3EQdNZr6/2m+sWgcYY04HNH24aDPV1ZT
xE/NbQEHMd16OBif8SKCEshiB1mm86r51rgNIsi8DqS4HvfJ4HrIYdaAXs/AyuBRibUJoAd3wVrd
CUUTkAo0oY3JoIGzREsoknP8hV+iNeFPwbW9J49Uw5KHE1yvhqqr4pBQSL5aWf24HdMXpAVh8anl
d8C9QgWJHbX6xRQsYVBNlzEBhVq0npsu4Ev/vgNmQGsWwOKTr8yw+WfqCv3K2XUeLNOqwuiuZtGS
45hFB7WRcvnwR5JSLfe7gadNh5e/JfWLzyzbJ2Hv1VfYaRXZk94E6Hn3oJ6eueiF3sXVssRV0+4I
bkOz46ogS3n1O6fAAm+dUoJQ1FNQi9RS6RrWG04NABuPJ+QZ5ewm4CIPyr+mBvKF83cqL8PVNxm2
rA4AGUTlonvC//xVyuS5jLrdgmW22yyQuOVuDKm6kP6pKWg26lAdLtaFL/z3LwiIDo5+Tbc7kLP0
ujJXQwFJntT4Ffuc7kMbzkrtS4XYl6+0v4M7lzh4/Amby4LWStnXSTSuHd3ESdC4y67CMDD/iIVq
tGMzUNVLvqRV+qJufqTJb5pG6nU4Kz9xTZqxDWAuy5ebRQAul9TEIrueQwfu28wYuoYqwL15fM+H
GtMG9vpOWFNc7VrjDTSWht+r7/gg8OdNDaiTU+axMbCLvaia+SXWOdnqPgruwBU9XufeMwRF08ef
34WaSoYNOX7ffIY+HoBov84tA5LArXi6g+TDFDQu6WsktJM5DKynnCYgUlwITE8foUdK9W4rEheL
eUpGxyYotn2rofVdHH9dKjtE+owpwv9kHbRlY6lle40IxIFPleXvRfdb1QEQpUH+hLqp+n5lJHUS
GjqTQbHRDOhl/iKKToxbQr5RUVQHJ4friooFit5/IfYT8EwNbn0Iclw/rx+uqOhJinj4qaxLyvjV
lwj3vsBP1PR5OSM7PXnl8pnTnQ7hzeZVenF9v9BmV9p4GWid1z2mPp4Tfyaf1MYnhwc5AzDgTQyG
X8iREuE6K2I6zO0r2bNW+CgE7a7zY5V0YGewyWhR8KHMD8IqvFHAQLyjJZGRb0jPYXcWVpEf38en
CEeJ75pE2PD4KjIdxs7PLTFwvf9wDO8wEtsiUCYeB/DS0QVnGwt3YQDGBrzOz/VojD1i4Qzg7yeR
DS9DmjtxE7Bkp8zKABBYcHfcBZMXilft9JTMPVAqaqX7vbhgwSrC3wnt5m0X5BABy+ixvixYj8Tx
VKEl1VldLyye18oR/n3pgZCZ+HzXej7UX6FybRq0krxAlD+4ONNLREuQsgvzP9o+mSVldorEa79y
HMlnkBmngL+nlDXTbCxMtaJP9yAOYsYUOt//1VdrNnQ9TS9yDVMELJqwkzhXlHUHjGqbMeJCf4MU
Dx4J9xp1JQdJc3q3TiyF0eqEo3QTiSwQU8sVIEaoTglIiIBhm/OKrd2lPW5REJwQRrrnfRweLR8e
QZANkJlykr8JdMNL1XG18VtFFSKn9Owqxej2/nnXigVTNl5npy2uj8UFef70bOZb+EfcxKvvxku7
tEWhko59T05vRpG13c2APEenkVpLp0oBAZpWfXoePpJTO7O1rBCVTlSvx/n1DASMFAoadpY8/eUg
SlTAtMJ3UJHhSA4OiIf5wacPdqO39Ph2WYufTgvJFpcW4x9iJI3eE9BGfteCmZ4L0jucDVHFY/5D
UixoSc6YJZTkw4iS4BdLsDrp3DYuU7ZOa9ec+7TzhOi6NWYIidETjuYiZegEOQcJT8HZmjy65BpH
mAvCiKqC56Z5WE5ag7rkd10YeJn5Vgo4c3GSbl2GlnOVhCfRh5lDVv/n7D+El5LlYTik2Ug3ehis
uPnOgws3RA+IqkuwvQ7PeQyChh+An4uEoIaJWaMhOTtpST6Z2ID3L1EaE6M0BkD3xGCGSTYisTqy
3Wch4j6Rr58C6Fgrt8Ema87bUZwSJ6lUR/yn59NRVd79yL5uZcAi7dAQd/3yPhU8nmFzMYkqvu4U
nhQ4Osn3/CmeOpma2eYKFfAkZjxviAwHOSZLqRoK1CVFRmm3mqNZRnqTNruqVTIBueKC2sKoHKul
jv/+/UK3szwj3MynFLYMpYfam5LiOcGQCFK0PZfxSHFmmgsNU8wstTPEu+KbTP0IazlAy2OxPM09
+B1secPq5LuG2ak7Fwu4SYWVQ/UgFWA8TFRYEOZ2hlzhF+esVE/7fcQWLkjrRjYFG2YvagHcUoiq
YHFB1US4pp3vO9HrLsRMM1kdTtCpSxwzk2SPrcqWCZnb3OPeyYub+QYaBfezFr34qzXQBEfFglSO
uhuk4ekW9yIgx8hNfGMYaPKSY/ygC+vMu2MyTMoI/TkR6gHUQh2y9/pjgVPuTxbGbPQCarFszU48
MbT3Nj3amLusuMCnseO71PEfm2v/vnQMjmnOO6g9DMxQTsb8mryU2YrMTkJ4iWJIm3TF9q3fuBxl
GuJF15c0OUj6REW4XtDvnAgAHjjFtIxb0XlesTy2mL5ZMit1DKMwwcU/T8pHbTXo5uZSaXczQ+JT
hDFXXJuehe2GrghL4QDYd1ZgR+WCbVVmb1M9881y1jOyP/vFm0NIrDFNHRmT7XSIIrV7AB3QXnJ4
047j84wvnB3LUgCNlSEk92w9Dj9lvaQicK4CWcVm64wrdG/GgIyU8nse8+cAoZdscWN3bIg+SxTm
UBMafwisY7JG/WVgsXOM1L1040hnyJO7W7t2HwK0SZoeR7RT8o3Tmoi6mXH3WCkDjayj9GyNrIuL
+nzLD2QdT79zXREF/+nOyZHJps/03loSlJrZ5OJ+2UlFG6t/bR2y+LSGHEQJKnAs/kKqI5GBGPJF
pL0jCal7LqXggV19ADQvmUE+PAy9Q+q64iNaROKF9XhOeSWpzmLWamsY5sZKQVOWoS75PjTb5lNb
C0kogGZmoGklyJhKMFIYTCGlWVMeFyJ5gakqXo5NJCA3eVLa+hw9R1j+5t+4GSvUTS78Uo/GFkN3
A8CVAdi0NqfKpJxiUjvlbAbZaQXhLZGkpx6Pa4rOhfEivyhrVid1Oj/+sRV0Sw7Upuu7k/WDoL0Z
eHI9+6X6js33AWmcLaWlCdV+nHNYA+XUXhjqn/Zdo4oStgNI0Aa7LKQw/tCpQLOPookZJhquRlr4
ZI2vMuKcSL0XQkD4RUs+kXSmCp33JpPAuXfDjxQpsFR2zHXox0EeGkaV6mXtp0ap3L9xkIRFGl7w
CJz3YME/9KpfasNOzFEckNwi/XIT56c/biifWlsZZ3uraqot92hPGWT5w5zMZPWq7ieLKEGJ1BNo
OrlSjkuCz6E8Dq4H3bZN51dM+gQI1QDePBgKxreGnmsDBKJrrp0XZk9dOnADaX6uTR6/Wmvj8HbZ
jxvPd2YCt5JaYBTm25OL/Z+fGaqsRcCGOomc6fHPGcOL4KU+tW9fhdDwCjF6dpiAMNOnXLYAIeTs
3wCH3C/2Y9NNqpXB0sQISSJmLgtwQf7bhXgXxnlYto2U25v13JN97pnpRmiM0kgOjfPIa46ElVWj
GRhYP0GVFk8Ok9fuu7fnjbGTKKIwiAg1TJNOhJTwyM78mZjbTVqnTYtN3i2krkTseEqoUnPMSoIW
AudYgcQAskUCP0xWMIaAs4cNDFgXZa8+myLW/9LwF0gLuBQGVt3sH32nw/9cHO9d27Xom6e8oqwT
bVDDqPlKmGSVtzpJwzODAX4nRtTaJbxBxMs8s0sA+tnFnqz6Gk6p5awZ3pjXBm8ihVXMWxnEafIU
jWpq4kImnfRKJtCknqF9yYTfK/+CjJGgvtZRMSkMGhFzK/oJ4iag1b3ZC0h9cKb04XrIK6sXg5Ec
4ivyr3k86+9AeFx/jw/OXm6OmmOdKDOZ6L7h7zuRFC1vGloSFnaGNtLddsEZQhMTi9C/GWInrhTI
KC79Zhs/yTOtYmMJckjH1iOWWc24Mpg0A0WXD6sC7gzrqWAq0iZ28HqIgkYOLBLC2I81eY5NBPtp
/QAdKyUy3RoMOLFtkNQ9Z1XuHw7ococENj/XDvq93I9oRtc1JjOuECHoHIjBUF5S8Iptnce8ow5K
2gQ2hlIbXNn/B3gk1ASuyO/UggvUCDSuH/Nd3e/HVyP0OW0NnlB3Fml5WtHo87Wg8GmBXJL2Dexu
eXQTAw5O7NpopssSQSCP619PiNgiwCiHfkguXZDuj8WMAf/pCyDySdbzPDCIUv4sFHrB/EyJuKJE
4naumX3m/g3spS4/CTGTixUoa+nCTeQaOrzXpKnuU6xPTfd7G1yEdeRk4eqVVs8VVBzSQgK1fRl4
fd4DowrEcR5pxbHvdNonjulE+aN7oXw8+DILuH8NMAyOz/5JOkYxJovRwfT7WyUsb5DshyAeyODr
LENOM/veuOi5DuVf9o4MSCNN1gS5LIgFsOOtRWcAUih94F5K6XF6YSp/t7oPCJdbD7uDWEaGNXaM
AZJXvIxaYydsCW8qvaAkckwbEeLsSY+1TVYHyv3ZOZt7400yH9FSWks+AWcOPKQFO92VtgaqXJzz
FvSFERlKsyRr8EQRBBnl4wRhEBr6hQu5ks1V/mDvIIE5RhfJdkewL9IUSL7tqZjHCbKELiFmeNbb
WA74yAUAFMgt6tFq3MHlhw3M6T9sRUSNkGMF3wv7r+oMZ0k8OwQuOxBOByfGFD6tsRXYWYbqMWB5
D9E1WmmdIfnAKA/bdrqHcXSv6OERhslcrmJZ3sudolQBCIWZ+zztTwV+vhMtCr1sY4JrIwpuH8e/
nB2v7LVdTRHspb1OkcweWoM234diGuDvkceHwbA6dFKnIDvZIzNMIBEypy2VqQhL8zukg2iXGD17
RgnbSzKGztpm6tGNCa5h70CUY4mywYKV1F7QF9569NV1q/8gbQ/HNP22QABhRWiUJQtAHvEKisZm
6TaxM+s1iAdMZCnV2G4HEKunckG0QfTdLoegfzbzNNNZcjqQC74fdpoCFE5TB7bexnLu+oobXhRT
/NjjMp2+6s6wgUunmu8y/IK4DKeLHXca/618z1Bcqk5xeZVdCyExp37yoz+s7ieP52gZdsJ5E1Gt
lcGpV/0PBO/HRicExoFUfXhL5w581K3W8ajMqdb+aoFY3w6hiWZhgQ9chIsUA4s0GgFGiu9V6Lwm
H0XCVi40Ldwy6M11rJOXHzTXfixJXhUc8UKvhylFy+vM2wMqMU3nEiOxiFqniOZ1A8RFdmHDcjj1
/5vQbwY9f3s1z7QHp4tm8gi4peLSwumgRqaiYTwSWxQlaxTV0NtWK5R3NgSuJ6Dm6ev5mQ7bnR+O
XdzeI55dixx4/vufrIkx3l/ASW7EnI//bWWEkIm2hszOjjX2amh0FjjxoO6TA1qDYWoGse4K+Tlf
5Isx/iKPsJr5/YX3DTDeVlT2Imi4QBnnU9nOBdjxLDcp/epkpWQKbusynttfbYMPaMC+x8cCd8r9
1x7EaammDP1Gi3mHVTkAbBU2MMPho6S4VqM/CGosrZ4n2V/5a7RpBhCgm3VXxxk3K4u5z3eaV9yj
039Ey2iqJ7ZugzuhGq34O/BC6Lldt3mtywQr2MzVOyinRgJV5z3lw/yG0PUhRnV8biZFKGyOzdOf
f/ffxlUUrC9P2tWdDDazKUrPQ0Kk2dFJQPAe0+I3msXFjC+qnqeXv2jHYxHFyJOJlyKG3BA14AbC
L53cIPbDem/x/1gFacywZGGt9/Zv6CPAv1bogqyoimYHS7A3eMsWApukDv1JJCMq+K4s9Cf1LKGe
ZIIjh7O4ofsvd/Qk7eUjCMMO+EcZwx2Ph37ZezGSK3GvH/k4cjwp9LWhVexNRkWqsbTQ3PRRKqPR
k+plkxVzP3W2f7hGT+/+aDBxBHyAmfyi8uAKUfJi9su+AfIccthizy87c7/6puqubBkh6LtKrmoT
8lzciMdYXNInt3yrmJ9VDbuNILaCPFhSmyJK0A0M3SWBfZJmJAdI/MMr0p8EUMDzJ1zdJdlbxzhb
1nocWevqW54TtYP9VBi/DampOQ8Bwf3jO9sL/WqWvbpSwbw90wJD3syRbEZcqfJcUSCXBo11XTLf
o3oiticSMUpPEWEOHqBnsMbwj4H8tiG0ROLoycxM+dYoL8Rpt5qcGEbY/ySFkvrsFmHeiMuDNcA4
xgLMhBFhmKrOL9a1YSHWYp5icUWYSsZPqhjrPdVVoC2k4q8mQgHjbUHjKMC8me/LU1Y3beufUd8G
HSGoOBeBVZuOJZmO5vuew4RaQNRXmx/OtX5o3xZq2yK83ltQX3JCiMJjWSH0lTEjH+qX6p4Zhl7G
vPXMmCwxWlOWpy5CODxqhmJZRdlvsQFaxECHJMrKy6UHwe/LOnytmRSmAYP8pIwt5abP3UC0n71E
dDXH7FvlyK8KP/QxdAzBTiPcU8wC2cRY2j9nJRtbXLselo/OMp8G/tJKBnv+4jE6oyOStkLxlNvE
P47wwmqTpBi/DAeFRvUxoqu/V0+Uzqx4yIJR311he3Dve/jGSRCbzYR4Yadczc6JC5OCiWYhaYGb
O7JcUX/wKFDMzrINjMz87Bk61iSnEn4BDLxQNXVu2rBq+J6UjsP6ToBH573xGSERCKX8hzmCOue4
6ft+G/cnSVCfazGj/9y64uiKv+gsKFzcCAGjeJygkbqLbsEIosIgs1gUn0AZfNdv0JMf1lDdQWuK
JIk9meJ/QWx5Q6BbAQKs3VJZmKR0zmtW3uk4eZXcNI3m/HubIuF7k9tC07s/bHyRPu/ths3ALexA
yVKJXCwHo7IgaUT5ZnvUi2yBDEphvtjRGp1nVQ1oQyAJmT7iXSMCyYsNx+/LEEBZ5ocfRoPS7PvS
rPhwgSfJZCNyqlSCXYboMlnIZmbm5lVR+XcB1ExQOVY8MZPrcRSMCOAkNnKJIiX+D1sHM2y892EM
RE44zPoofzMVmil+x6zlQ4u0oKJ3Zqua3uRZ5R5OSR/ex5RJHdyKvm65/QQMRlcVIuby64q+e7ca
9qjUltoP8g8gFqO1k++vXSuHGVJdQzZMLEOIpMXgXwA15t9BEmWJmGrx0JczGdlnXWAXBoXbdml3
nh0TN2pBbmyFWzjww6NSkitt16Zt+NXLkaVeNpUDXYOC6RP9Z0XxjDu0ID9HOW4H5vSEEvW3o+5k
5OpfEUUTDiHdrEWpunzz33ux+N4/nkTsmm2zAQuaRtCmI7MSjXcLGy16J1FPSjzyjXJ9vT3hzOZe
LLjIkMQUYNArhxyLaq6F8ekv9mJ5Drkq11CyELi+U6zfaQbXTRWquMphtm3+wdmo7aKjYXYT2BZk
WGRdUIzCMyNFligodkD7vLGGRWRvzylutdx7wLM09pjNs1FuYgi38pVFMpZhpciZODhtOj0uC563
FZeeqQPuUlpLTD9CNX44QSXH1nwkBpORPqEADQkroG0AlEmoz6cOMpVxXn+glArpB40ikzi5yH3f
z/EOrOXk6wduvqBu7N5bVTGdb38PqJkA7aR9U5ZPEIczQt5ow/aGQpQZS3vZxMRELfvW8MbDcRt5
Kv35odaRBXCsDKPF2DrKoPTZDOEtTUoFYfagdx3T1f+0rU+og8qht8ZH+/QfIMEsI8iUNPz0YLfx
VqoQR1uiaDvUY0a1uNcR77Il2Y0WMDdczeU+dLh31bA/1AZ3cP5zoeZisg2Kgs7Z2OxnEUC1da9Q
NRVixD6DRuB1FmuotnDnlnsMhp8np+eBe6P4iLO3Qd+rbgGkrWnxzfbXxRNCuO1vgGlom5Kd89T7
diTqOpCH6nL1PMkcUS/UrUpHzVGxKzie2wG+YTs6a8Q8ekyh1DS2yX7e1Zxy28gCV+tK6ESQEWdm
4V/cgEQmPeRPc370ptxwzros1T6qSpzDMf1Y/coYPI4+0YVH+BhamcsGTmd97ZvrkTyPxJmNdfta
t2ISLht9oHIEHeGkPk61KJ2IFhMadcCa4r6gp960sWK4HfK183ZPFRXYH9M8SBBJhZ+GwR0UZjnh
JVlB2b9tc1ccezaGLu1rc4mCRZRSBRAHkGftDnxrBNfUUJJ1APivdWfv4eaRBIiXUmpZvrJqO3Qz
hJmbEakun0vinD4liKKaz/Qkc49aZvzFHdv0mxy+1uUncJW5pO+JJ/PFnrnnE8I7d+mxPh0o/rSL
pI19kdG1baJOwxYQvfySDtMQsbTiqFF7ozP9+oI/2d0ugyDX0ZWcxG4f8oitpvYkd+sYC97gdJNH
70nnnCdtzamsKxn1mAZYE8Yq/HLtPYyg6tQeYAJr7h4BvTAu/uexPaZPA5jSbzzoyt8HINFJbDci
NP5DupUnqunS1SyohvKSCNrlHge0k2SVcSDZoiZC9blWdyg5y6j62QTUdtHm+Wd850fOmqEeo/wI
Pj0nrBpfxNh6dGBy2GcQV+vKjVR/sEeRi3b16A93RAzWhdTdiZcy6GmDw6OULfU/o9O/kTKXISbB
m0d7cllWbzab6ywiAHOLZ9jEBDbXyoC108FZ4wYoFsB+Fj57qmkiUXsoGH7VYPiOqps1Z+N4Gn6Z
zbkC8vC5SSbqEW/DhmCbGLQbIiBpCobCbC6prCgx76RpaZeKsEYsMM4sY0EcJrMyVqStjuNgcvEK
k4MbZ1eHsR/eK+UoBxdH9sED6bMRGGNmbbTyTh0MmEtzWjMwaf2PrfFD+ALq7Z3R5VU9N5u/B14J
S/wFG0gOgCB3avjwIch09R0hU2rlWG0SZZi/XYYJ/A7bvjlg05ASg6BLd460XwhlhRcFcbZE6rx4
mOpjQ2pD2gm5R8Q6YRYNP9xAxHKpHIPc68m8N023z0TY91+GO7/QruKPcSPdrTrTeXLcGFoqJWjN
nZSK0O4qcHGC6KPEYJ3zWtCU4AHyd2/RW/1D/9tg9KDWGIp/jEi/MtUeTUC6fcDlAklS0ACuiat2
LEKpHLca2bYNtil9lltDaN0ZM8PNgVr0oCG3c4NXj8s1W4+Q/imH38J7jjVEBiFhW1cfvZ7uh8tG
YAxYStYGHKt9yPAuQlHVAx6dQdMAVgYreHv5SbGMogHzzBr8f0twM4mzz1oZohMWBliBlqiPcl7q
oZQ8A9V/zqvlyLsLui17TuDEtQVc7XE7I6M5jJpghvHWKWW+MkxX7vkXWshf51Ex7bd0E6vw3t6A
atQaM5OPeXwHvvTil0/wxRXj7Z4NkUjwrw3vNom9cnW6FoZ4DGGjcDc/QCLGnkSdC3dl4AV0amlj
EyVfndLoxiDy4A1z48q/rtr9OEMQirvuEtrqmiJnNHpoQg1J+exMKUwjm94bW9WKyizS3YUyUbsJ
ILLr5WOHul51jLlax6QAQoTgSP9RWlsKawTxS/DpBAMSpZxkGhUcEvM06Xh4nFP2XpUIaSeabekL
ZfobLnO9LbHFdRGimmHiqvbia0/r7MCpbdS0Voah/07oCjJztpMEEzZTPPZ49ylpp84nF+855bo6
Dbyi4WJEPzWjSgMNBc3Kcul3seNGfYHDioKcfZTOSz5RaVqdFwTIKMCQWtNPc8vpC/7R09/PRmnT
aLbW4GnEHnTgNQ8sF6F0m9uCIgCLqB0rMAvg5zutC6xZ0FxK0wTfYay9YYXBbTiEKO+FQgLap6aB
ctyNFlmAIio96mwscjxemlCtSsqCv9PWTQ4BkRkYfl8yU3R1ZeRmzbGjbZHdSkkUI7S7VeiDWcAW
jNJi6pRLDAKh+LnQPKfNwEJ3B3FoVoUk32sQcsyXa7SOkjzPIOh6YDAVnPAXLZNZ7gtW4GEOpROa
59C9TniuJtKE9H7CfIBwUah388qTECMpHl8OGtNXISIh1Bv0SvD9kea+3beoHLUE1gQPoMdLxbtO
uuMgigsEJ5UTXfhta/nPmTLLwB075cAjkC+MfRlscx8lg4ngWQljVQxpcsBUPWYlxHn4DMOI5kul
thv/IFgb8pLcL38kObz6TT11XExpX3wG259/qftzret5oqQku1ATRzBMVWR2H2cVJalF3b2ZO9Hx
B/LcHglX3SFDsFNIwrYWCzcwCqL/d78qL8Tb4wFsdr57jVNWC2oYr6EFDfeeiUvhnAKXoj/89qdD
gISZTDapWEyJnrVfwHsWGtVvVfPCkQqnJ5H9uPcvZ2F7FovrTiui2tZ5xUnnWsEM6dG4o4JOKcxe
C3Oh8EXKVPOiZgocRIhTnQmyqtxUeujv1w4/985rqi/Lii++gBDzK+J0GjjkwIWQtu3tegtuxwTj
8Q0JnTIlkca6WZiMuXRJ4WvE/h55fWwi6U32/Ttj7jsNyzc7qhYt7NHYl0nx20VAnV8cKmtJMvL/
36IbNBFss2CgbFzeleusfWwzAFzeiQeg/IcPArgTpepHFsMabo5adkCyrecGbr5/dpoR3yDi2twG
mZq3s8DpBLk4P3Z+fzq1MPSLwAcC226FUtD6kmiXIGA+8lMPOfRVTAXuDOltpMBleuZpmrMeDnKc
VsNOR6D8OAuKmMFprBMrcuyWvesZqYBVzjEIgQhdoYFnssWfkisF9SP4uCdrC7fxPf9F3TcsCs6K
RWOrqfvWcSBgnTi7kJroZSFyho8ayPHA1XKjMKfhtQ29dKu+QYGBVtPL9LaVsmcBOgrjf0vO42+/
a61MAikwcr0tzPeUefIWZF1E4gOjXagktx9nPTLD44cP2s8dPw0wz+Ma3KJVFcEne9pZAHyCpGM7
qJsQTd2BzZucq9/ZJshhaFgSISc/Q0dDECpfipWmIQgej3VZFQKvKldXWBSIeRU54kkL99B6/rhP
JAyWEbefOylCeSu+sXc7utw+oeo5iCVW0Ny6OwSDE+amvVRZNQ8/FhXFb9V28kaPdOq339oPXB3P
oH1dN+vAFmUMDNrJXw1u15eJJH0k81kyuwJBR6ze2mjOOTy1uBak6Ti157tjPdX4Jtza5Rp8E147
o6B+Iv/6mz/TkXAq3ie4K9H83a3XbDtYLwWJnV9ES8+aABhmkPR/RAqGV3g0Zx+tFHbkcGl7HE/+
/vJDlkAhlme/nP0LYDfbNCjKENuc7JjzlI9Lup9R/cUp8YoP/8ShXpJqQEe+9nett5pCAdV4HT7A
deNPO98kLq+Q46MIv3ZPDY+/ObP+7OqvrAvbETjxFieLcWGV5YCbhOq6HdDUQNN/iH/gvgHiga6p
MUzJVcJk7s+Fj+zLfa59CPPjk5NFzNod18MvEOBErW0ppBHUU3ynYMjUMklCHNUd+1yjtSjI/nJq
d+bGUlLq+KenruUy7+4Q0GDIDa0tIwAKXRA1b3UNjzx6oxzSpEZQY59xdF7Q0jwtkWgVuUekum2f
e0X84S96WemEQosJRXTQ3zfpDptMXMuleoiCx1U0pOLZzKZvd7DcZEpY4UiQDCW3vbXpwHny021D
A6b283SWWLFEyfq1bMkZAasykYn1DkPOKmBGoLdv/FX1ZHm/9OiwWF0gmqIuIgjFECRjxqNWJyca
AGR2jKLnof9Ju8EvyHSt3bEER2n7KwU/eNochyu1ps9xuZ3Fh6RGBnndfiSX/CtCPVYlf13feHCu
HSzLpjGRmSTqMkBbqxySpwJwTaXUoecKWbPgWY23wpzED2uQrrwDHJQhiG0nl+cz9JWPkiEdgwnK
bSYQ1qkayqQDT+2IHl7aV/2fLx6Y//wIBKsXzgVSNqllHiIuo6RdHB5456IJAfHeVV2Luu+eWgIq
Fh/+r6L4am9tzDr3FmrK6astP0fKKqqQVo/7qUA0Z93JvrfUNu5QLsl941EZoxPmv8+lUjVwoGmQ
T+d0J4MNBzPmeFFft05hpjlkKJ0YpiJqmK0I0b9R8898WRnzDExPdzgdccjtfPSyfIVr98ujVUow
2jB6UgbkDSaVuYB/ZTuvb7CGSSiSd1wi0D8vKaweKXqH/vY1XoggdDBWCdgbIsSnkuYM4SXr6ZcM
UIQd6q1Zl2tOHAcDaYzWa0tf5rsyAjD/THho868rcnU9l+b/jTAchdGgYEKU+t81gUpZvaLWqcy0
XUUX73665BUvwgqVwdCLOItZInWSswL6Ddhn76wbkKv5/TNetqG3MHuxMuUgg88SxtEKvozsm+Hz
HLNNXHtIm5xMI6NlmK134U9jB/ByaOOQvByv239YKlTfiHECweAPIra5pnHhJOmxitJrUpTNzqMu
kdXzeTDT4Mv6dr4VGpMfr9V8EG75KYVls50yQtx+iQiUMj7jdNuQxlv5UryimcXnMypmFLufhzIy
UVi+/+aE8Zl2vyXvy5TrgW+H7HzNYpMrG9VhAWNquxPLfHFzOmy9uZP0KkCJ3M1UR74NWe9c+ORo
iS72Bv8mqhNHwU2j5RS0f5xw4keeK7ILNjeu3T08ZVRs1lDX9cUH+yCsbh2IT7rQFkq8WFdxeAwH
hzV7RwJtFW7oi0J4LwdY4bfeSIO/XcnLmHzoBB8hlwxnh7AzmaT90Nb9KrstelOwpqGpMOzWU7u9
4aOn0dWbB1G3qaHwXoAGemUe+wdc89lquBQBuEcCNX5lt12Bl5kHrlwmSeL5d3RvdIWTmcv6CKZ/
0DounpEXIgNW2RsywUOeIesLmT9NJNlf3MTS1VAN2/QeDVLHTnYFjAzRtAe5U4o+suukq/cKGFHB
70uH6A3yK9RfHrbqxLocaWMQuUgPz8uPhm1s49AikputVTVqWxRMw0DonSwjPI2yE/iflaHcHS6f
1HGDkghPGtDCZv4504Ks7DqVu5UzULIarKiwuzMdJ+hHFY9ffP675/xvhgpDdkoHR0h+/srKjbO0
0LOHMLiCFb14gMO2hhgwh62Nq0Za8B3UQn90WXQzoya/Q91oTnitHhPWDrOeQlqFbNn1qTUZzBlA
VOtA3m2+07rprCTTtuwFt7A+ObKAHZrf2xVMOt6YjHDeQpT/DTHkIBEmSQUX5JmL1CuEMdXc1PWf
T01zjUePgglJRAkQEmHziX7VlhtVDdfL+TvBnt4U5UUo6IT/LgEtXgh6AbSbewwR1O8Yqd3onSnQ
tDI92BgjfNF6Abqn+voPyROTTEcMcRDZ1F+4HYn1ue61s/BenrOx1gcJ2VLG7Dk3d90fBQ1CzAGi
zyOkIdLLVDMSL/5tbJyjoTZ6StbWIti1VaAlU0BRPBLgta8IV2OrC1TPtqJUZjTmQcfoUrXsbi7H
QW2CfXj0d/o3/1qqCmulvT0LDmcILcoBPEbdqJ4/dBeTGQ/A497eZPDAIpnO0tinfILzgKc+7k/0
LvtO/BZmMu3Pb2yvMxNyS8D4AiWtlVmqysfn2VXJTYTBzEWCIgbUXuCDUUbGxVHBuEZyrO3VJIKL
Di59Pbpvd0za45R/fuX0OG8v/lCFlgesLDd+pZw1IZ4DAh7hjGJ3E5BjBck0+JrXh/lsrT8gKgOT
4yhmFxWWEXdryPe3SHYWa3J8OwuJWoQqqi71VC715GuHVbCgx1eAG92qEpvySkrDNreSBHfwLP9Q
VK+S0Dmz6PGFc+ZUanjSGfQSl+mBxMraRUjQTfh4MnKNPgA+FSsIvXGhmbarRYfsiQU74Wz4zflW
IzpD+aZHS9gcsDQrwp9Xc7+95PE0Sa8p7imThn5peSNe6Zv1kXmtQ5Y4zopkPR6UWCrXgKU0GId7
29H3R3AGXXh07Jp6qKL3PoL6i8FkZ88yaVJgB+psUKDTwOoUo1zCNOup/RfV6ejH5neTZ1CBRfLz
jrl0pt76ULhCdY2/F5W6cEZPYSuHJcxNm+uV1JKmDmp0eW+QTbFEgoBoVIVaYYg2ZYjp6WxaoqFR
cLN1LNJlvmCoPh+v9kvVw0iHcZKQoTv6N7UwydI7m5nZcAJCjFEcNySudAHl0p82NLhEL6Lt0SSN
Zhq/ids8MSny41x6sF+bv+CAs8HCBrPD/YkjoqBgHqA/FTXZDQViE4ncNKOFvmSna9HhF0+KuuED
oDevcuDAwa20YcJfm4dwOUqjZXI2bhyEqmEhTKIU8OAfrW+2YsAkKFpZi+RDxs2gHud2jHRZ0hAE
nMR3IKll6C3GsPMgnPIaoapiUTVwz++ZiBGesk1dIbMgaMc3fvEy339ntqJd2ONuUe2m7AHJq3gD
eMhltkdwLaT9xGsYUwuCsRRIj6n7TDIYCfvzpoKGHFXyBgsKue0/LWY0STFi6p3kVAwWUQOIt2zV
AL8g0K/dmrcu9gq/uQ/pL+WyjPJpUf/2TJoSJF7JeOVoupXG4dht4BtOAOHI0epqVxuYFLuyLmii
y5AIMMdf8XnNVN2LAW2rxtjv47J2XERyZiE7El1wP8D5cipSRZF5CYQsHKk2RKAmLOrpd/9nHBLa
NtJxDdusRhhZVScCORus+rdae9Fg96ff7khKVw15CSIB7Gcb8kc+OnFOi6qZkaCvaWY2yOwYBsps
l46v48YtfalNNSlh1gzJQeaJB3YVmlXnWXVtDVWoTK01j//P/9vMz6oBbPNloAhnznvFUixez62e
DypKXX1SVj6LNryGPlJJSJU3Zh1CWnFx/cyerivBPeAWInmHmT40W6NUJs/uIoWqnUK/M4cpjKB6
gStp7HJJTJhJp/aLO2n1KmzKjuIpUJxCBkoz6gUvOnF7Rs36goF7cEieNhI5E3z30e2jkaVe6lak
OGa0om6kMvmAgzquQOalmJtTfeeaFa+OgjD18A9gMpbb+YIxmoyjP+NR4EMCQxMS4PeJuwcQ3Bpu
LQRCmz54O6FPSIJdaTtdoHNsUzZGTDCfyfaeH6WAE6p+JA7weA6whKWlCItdUFhCYMI7i/Sh3C6J
0iN7PSv8juRF2FI9/rUi/hbQKkSNdGuO8F7Hno+WgvRaxHlcG9/36WPHt1B+qbc1ojyDEilm3ESm
xg4taedyy5p22rq1HiH21Q7F6CQ7Ix7xnyVbc9uTooU+VRuTne3PISdo1lTv8hcnZTvjnyTg4bQN
4RyP77+9tRwYo8YQU/CkI3x5sPraPlXsqZLzeRiSxJ4hHRZQcmRXeIdUFRF8YX/oYsOB0eh/RR0Q
asQo8KI0MiBPEBjpvWyR3a/7b70ingQlsWYRghICjAKLRxgadHxKdpZoP1vSn3h1AhumsbmDFc9H
eXcM/jIJyrwUovJkL3nR7U7HbQ8Pwc45LizzQXVLCeIgmdqrKXE1pNhmy/tTON5rarAsQ2LNaZFW
ap0j7Hkb0zwL4ex0Re+sdLN2lDLbL6rkeI1mT2oq4ei8wVhHE7ckpxvCg28Eq7oZSvYSJK8+fvAm
KCFP2kgSwfkK+7YQa0DMFrLWmSCmCdGl5QwiK6ni7Fwe1co5/YgzYjb3yFSy9mX6k8mjYXOkqAoN
ah2zjh+AGqdtI/rv+HCPl99idjMgtrnDYVXwi5bldEqJsKoO+Kb8Q3+az9Ji/iqKb6jJI2NPW9za
Rf7k5m6SRflyfUXz0Iv6lSEIBHHsj56V1k/Qkp5hVaDRt+X0aA+FTnIlZVttKhuT0PaC2y3KDuH1
qJR7Saa9Wyet99cPV7d0wC/opBsCEEbH+ymT/8/A9h5M5ttNgQJ9UJglieda7GOpVdPzLmAKQLfB
D3sCLp523IPVZHn291zFUFpQE+oIhGidpVssaW2/0xHFXnD5pIdiWkegi1qS7w5hkyDD5BOlWspZ
T+K2xIm/qvpHb3YUt6MASF8cBj7MdbAoIsJJZ4b5T5vqX2oo8iOtzcQk6NcLZNL5KMGRtLxHrnIn
uE68N0ja2xcTjVu2GhV6cQWnNR9vxXnUB1ZdGeWVfzkYyPtZMQMmSJjG6uxv3FC41zsbPly20bGB
qpJN8juqkMhehUGolPXKXgJdzwUbrPwJ8rx7mB5b/hxs5DkgODo7sTiV29q0gVdz7lx7t1k/BGRs
ho5Y5gv0Zj0WbaRKcXhJih2fO7Jln4OhqCTi3HgXHfhRANlCa7RX2BeKOEjBjMxJYSQ9O6OPikub
a/u77M+uL6mgN8VZ4UyK6zit/Ir5wHh3QsOq/C27pHt/XHv4HUvXAzGtV93fJYtFU0cmeh4gDKWW
Yve0JDiCbT6C/nba7FvwrEmhJgG0L3SQy+B/RGWehKfIVDTkI9m7JPxCY3Wed/8SgtsLwBAUloqk
Lc1RJMWyHXz4XhQ+Ne5idP3yL5Sr4/R0Sk2KOKgxMDsby97DUPbq0Yz14do658J+MeAuh+bEuL5x
qyft2763QL24211zTPpCxoT2LztI3N+ZLOVnkPRYaZ7ON9t7lMRJgcQf6G1A9weKcIUI+hXiF6FJ
BwA0hUIeZshtTro/aU4AKxk5gUUtDDnwAsH6h+7hp+B6RWEyp7n6ihchdPwaPcP3RBW0KOqiubrl
AvKv5qQkbAzaHmW+5MOvycom2J2Y1QYTdEU/GNyC7BDobmqKIvaRZri4uYLk5qVB26r4yDyC0Nz2
o8hFf4kynqNMrjLF71CTWymOzehQfUIcsOKBYNJf4k/oKjV4+fgUqSIhG2wUv7pAYPYUAMzFymr/
5Zx93gqWqp6ZFD2EfI6+bGShqVgDfm+hsRdD81AUSSJVbygIvyMzvQ1qjPvr6bldVPTHj5Q9bCtY
GidjMz0d9NtggS1xTU3syesiBSdm98ItuLYf8tXvAL4UtRyKBpe/Rk0WcTKr/8DI5kQOjCb5eygb
J94MY4OYu4Celd1H3m7pFdpXqo0L9U9BoqcTyiM8hoEgLb8CIOxt0ElPg0kalRrchVRgQqaqZrR/
zhCTkVP8Tn1XtESE3mo50G1qC/mRuYcTGNw19JD0k0dR/164C56DAUkJJYJKFaxB7SDyk7Icw3HJ
CYWgTQt6Gc2mx4d7b9Zy7hgQjUtr4X8/XH+JW7Y+m6PTn0r6DW5hM0lH7Ra+x3ToBNlDguiXSSEh
nU1E0dtKP6Zy9mYvmIt/V6YrdGc9A4Gu0GcWGPSqStiI1D9BjLifT8uSHvRVi0Auc0eNZHg2i8QM
MgsEHXtSqTB3FLGjIsLKfY6fZGQ0pjB8XFBOmFGRaaULuIDGeyRyQUem/X9nkndhyBhB47pnqCd9
sRTkkwWdNfFkdIhXTfwt2NlDEw0ICmLLN+KcNwFJUQFxCbFR2CzF+EQsntsBonwQUoNtVki7kuzn
B2+l90eWS5NIAPjtf9MnTDp+T0B1WMmxhuhURJMlbxzt0RJs0tZ1/sAIp17B6+zcYpEZ/f6ymjSZ
aO45LPU08n+FKaFG06sklnCpkKfWnk5vwmkMKRJV8W6zVT3W1CSj47rBYwKcgqq/9Izq+zPzMsM8
T/RC41cLUu36cp7Nw7CzMxh01qMWaqvSFxttzIm2gk8SW6FRMa71mXDHuSSRqpWBYiEThcMs1dmj
9Q+FwBdRUhTLs7wXmmTFgeoUblhOWS3a98+9g2Ude1WLuWmX5cEwcN6f2MqYCW1jSNu5J5WjpRIS
+oUuG84N3OmbqfzBcl3Cz/mZWXYXzE549cg5z90uqEQsZjg8vubMGHte0EYQ0j52ZS37t5LOv/Ee
iNohwRb/9ZPhBE5q8b9XzQ89bUDZfey1ZLd8Hw7FdkvzDKwaK0yZLLytrXIHxiXzPMN+PGy6Sl82
29xxUjQrcdyFt8BfcgDsFjJWFQBr+3R9VSPfBUqasrD6xm8/oo0PaoCs9N6HdTgzknKvK2F2pY9G
kQaesvJjeHQ2/KwGhp0cSqr7wyJvB4k55olr/k3oZ25J1y900YtmeWIVcThEXlKo5iYiUFfQeFfY
/J1QQIhrg0eqH+L1QFoDPBqnGMyW/f1w/kR5UYWKnXaJVgVaImM4DMSrJli9tQgN6UVnhHFQk5qm
wY9dvYi1xpotNvxrNdtJitjsvkxNLprH2Xa5lt+6W8I2+9Yq6PryycLcNS0flbg9Caqx2HcRwBMA
j6KtRc+AkwS+S2WrvawDPawH+Qp6vCz9TTeYvELjrTnxvTRz2jcnfTqND/LoJLU/+tIIRTWI22hd
eAFx0gxP+HY/BKS4jX9WsiyiShkCQzBY+MVOz5Ocfhisgff6GP9D4IZOy18OIvtMxHQ4mnVMZb0I
J4/gf5pJe0N1ugzE/g7V0QMxmm4JS4GM9ZkJ9iJE53r3ycNtGcj3KXIlLLZHqRUdy86ZCfZB3WoU
JJ3YfJADkch4flkhPtZWRjF5ffkEGphkMmKMx6RJV28WDUVqesbEA4Jzuw1mJoEmgM5mAaHK+nuC
owMxW1iHz1dPtMfFu/VOHFy0PvXzoW1n+Sm5nmbOT3Yaj3WdpaaeocYvJpZQrmM1Rj0st8XZlUtE
44uKJFc/M0nm4kCdsA0iFRqYQNT2DJw4Abv/A0rYpssgIXu1tZVkGHKvYpJ8wqhiZvYIUeRnQcD8
WqYFVT0wvuv25eoGuu4lxX2Z76M3Lp/IuMIi3dgh7VvNsj++wLciabotnpMLnjMuSnxI6RCHA8bW
UppwnW2OCN5PJis5Mjj9a8PKLkcO/xAD9Aedwgnh3srvhQSfbku2wqJjBcETJgV62xNBUe9h8Xf9
WK5VED/kuCTVE+7qy77CcoW16iS3sKH/IYrdUJ6MJcK0mhwiuBOhPpj+JtAIiu46ykRpvnGfTmdH
SGzHYchy3oiCGS0DmEhSeeVJGt5r7UKB9wmum1zWFoTNbOI22voYpPDAKr7BlhJOjIyniUxnNS4Z
uqRyPuvud7FoKywAxbh/TPK49IqjEUEuGfrivcyfE1xhbrmO5aFcBdUkeesoG2DwI2BD5b4+QHr6
HUeKrCt4ergleFPuO1bbhkxW0ZtxqC2T2Zs+zqsvDyKMVpiv/vNi/5yvp0evZwc0axJTFkTj4vFf
ipmvGfRYxWwBMYSRxJljM/iyBploUHP4fzJ43NBWoVaeZa6Sy3kIeFNmaMUt/ljSb4f4geC4v7tl
aliwb+a8eA617Nbi7FNO9dHkfctmeR+TZj5kuvf/jLlPOAWA12hPGrsehEP5CJ6R5UtcOrZZD1Qq
S04+zJYuQgaRPHgEtZtgmOhvyroRn9aIs8uL1N5EOZkbk9weq2DbUBew8I/yjXsc4dIQ2SG5Fihc
UD3Cfw7kxHDOB5E/AMNLIsxR/jUl8SXofAE6LIZQsJjUL9/6caxj2YUcYxrhEAT8C4/BBTWKLfxm
SnTPBICBFm5gO8szScpelWnHhqjMGCwABNgAyDJoJWYdaG1f7OrKrh5eWxyJBUc4pd9huFaN5C6w
dLXuNnEH9rdxgEVNNrLh7OVi88iIZJpfHa2yQAHwZnasws+0GT7Ukd78Q71g35VkefAtvST3P1X8
jykAeV952FD3fIz1Zz1qmz2gmUvI69aZTPIr/jp3BstApDCbLmhWjz6/PZnqUOQb47CMswT5apQK
uNMpjl1zwHchGs2J+EcHU6IhTHefPHnPF4DPVOBBtboH90tFsJFxEkY7ZOiqVlhBH+zoIAblEUFo
mncVtkZs/Ni+sykDMzKQ++1/XgKzgc+n+RyJZcXsDdoT6E5tJSPbFQiEVuMlLjKg2twvgd1fqzVP
Uzh8M+ZmXpHS6hs3qHPUQJV57hahCYfBJfCv3Oupnr5BXTs2M5RMfIdCm5doSCnLVm1JZEbS91wT
VCEJIH4KH5xQV+aMs8ND0Nn8O7dfA0+1AdECO3UCS/myPkNdg5szqqoA1u240XVcwNhijxPHA97b
ESbAy8dC1q2IEWjf9upMNjgnu/GBcrwSrsyCdORte0E69iEM3qo8UC9fihOwwX7WxtPyxOwtDP4B
fF2JyoKhbkqMhGowGsVFSrBWHT7loRW1iEzDEgoqpIZAco+/6Bb1vlaSRP6VzzO+cQdBctUH74Hi
3j/0ttUT6S70Wr0ynBz6Bl7w+c/GpPMzyXgb7lO+plBwRjMHPV7qApeaNrGdtDMfiRoBKAiDap67
7pRm1o+Bv53qqSH0COZ6ao3/5nz3irtyQWOC55YKFm9sYaBKfrR7gVm+jzlm7T+1ioWM7+ApAZtV
zEUGnq8aFdLURI5V6tDwlKWnlKQKwxlqamOs6g9VJW7Ckj1RZod0IqBybObxSNDBR6ufsQtxje+/
d6FdknI7LXxn6ODpyufk8b6bR3F1BEsgtohwY6O5R8UhZDjVZ1F9LeyZ3l1LvYn99q493O1qwN8o
pdgWSWdht8qPgZM7tkRQkSGDZqEROcuaISD9j9QIuUJBmXSEfxj7KR3e8TX0AUPcDiM66d6FbZqb
5NpTZDjSyouXGVFXRjLsEjsSLqiotypfJnPw2n+XUSHGHyrM0rdhKe8Chnop4C8sUQgdgJiT+Zcm
NgIsavS9W0ej57OADKlKI5+v4mHFuwv5tJzIYaoCeaOXcmeosp7iGm+nUBkbkifgN70NV4Ct7tc3
1Cru5A6EJ+EvHzEnt4OwBJJJh6/zLeQ/KyotKZHSOS8pnosucPRtravIq3lQNhUDhu71qjwVBlcj
NmbfSSOAwEhAHRNZu/MOjRaBStIAMi/GfFYBUohXWf9WRbinKLZG/Aj0WYqTZKBwjj5k6Zq1DgIw
worwcBlLhyg2//cAgoip65g3LUlZBr1Z3SAFNnNue7ZvROnoG92J7yfu8zWOLyE5tIsJCjbwARxm
A795vabrTuGzgrcKBd5TizKwx18a4jNxuqeOTbTX+mKfcuJ9SVEMEJQHhAqCH0fOMvCpzsjWJxBu
x9zaXmLVgp2ZMIGMv2ah+KjbU3FVZEDFnZ/y+9pdNF+bI/Lp0QgpxFNBjC8kCR7cS1QJdiKX7aMI
ZU9bUeDx/B0sc+bu+HYqyDcDrDFb2MS+kzGL23EA6vdoWl3Iodhkd2kvc0jiVLnMqyWT130MUl2F
3WTxOZcMNgS3EjfpPXtL68+WhM5inyQ+v/oVEE2yOcwY3VQ1OMjYWUlvLz9S3xdfVI8yQaZEfX5O
fWd4MXd/spWp+9foEHugvgl+QUG+CQpyle9+kSmDHKwILHATtut34UnOCDSQm26zRPIhL12ngfTT
cEhcb80gy96KXSdaGSDDRqQuWtWhTe0Vkueh3XXChHLf6JmGov8hjEPqCqzqq5Cb/DmueTg6TQc+
FFhJkmBLbFintITgFbzbO847Eoiz+HiuDHb4mWkQGEoff1ISmXnizR3zQtUeKr3MM1JJ0QwfSoKe
fRtsSTSGyZsIjLElzEnSTRhO1tbyIke/yUrxxODV2Yx8Y9Im2xwBiufPZvXJeuNRapSbKKg1nmb/
iGDDQTrKEXU6JOMQEzYTlbqCnGsG7z/cgzTPFskvqRUSLKmh0RS/MDa7PVgNmMRfwJb6aYljGS4v
kHllK4iYSFnWDR8qzpHaX0rsu43iltLuNoCyIAByctdtGHsm3hcPEpvL3ILvHec+u6hW5UZUidVE
0ymPfbzdKrZqICBA3ESu1IApzWIk/6jAL5gdueYuXrIxllVQY1pE3BhisyPhps4nEb+WrwMVbTDF
CodKQx6rwLCjdADZwhIzNH/9IkLShS7NksC18Uxqbd6JFEr80ey75MpMq6ufHzD0MUG2g2nHMdJT
vVRgJHDSZpyz4a0MQ19DihPm1T+KIfHeZX66knRWX+AcyAiXhV3nI8fyfs8Qw1pzFDAZ/dO1USW+
jGsenN2Epl5QKGGy8UfcRmmoMJV3P+SW9Zx0SGEqRYK5eLQhHr7WWcQAJ6QPZM8JEEfOoFFqDgDw
wg0YTJ2aqo0t1OeGsGvD2X+wAaw8zH7Htxo34Ho4H8Vafu9lh5/w0TrrlWjAKDB8eyXqcO7y8Pk1
d1E3poou831Wh4ouD+9fvWIC/joJ5/93ex7xe11c2+wptg/HILl+JfPr1xh03JYxJtJpdHECCJ6n
WLhJ4Zgu83HqrBHBvJX0kmm4ZpiGptEvAZnrfItWB+ceWhYXPEfXjm2osrzUGvChTzA9mQXx4scB
rwNZZpWLCnuXNR1ASp+pgleM8WXYiZdd4PYNEkyJigL9EQ3Lwjg+8SdJ3qCAyvFfkqWzvw63a89M
4vUUokeuz7D4GdVmUGOIkeCg22M5uq1HZxPdl+9UkOZEUnhfSvb5nxFrfq2K1Kk4PqNpICoe3Agf
vNQ/DClkyudIoYf99hF2rxA+UIyJNqBMkjtmR5KR5OC14l+hDAIAkFAkAA3MNjLRWDdDPkvMfP7q
wG+6H2mNfp7vm2bLAba3Bk0yb161gZbH6Z9/sY1CckGEXIq3S8MNEOG8frUhEcwuJNWbCJ6QpxFV
VLNfmt/iue7xk3JXkjYDwUD6Nt5yxf/aU/8ngS+W1YsBG2iAqwDw+/g79o/mlH7I4IvVG18qC9CX
1+wBtc+Ia0p+3QGXU/m/zRIFu7KlV8HE6u8FuGsflPxZQY8Fom+JY7Pz3dvK5oY+/Dn+YyBUOurZ
kENeo4H6spEsruXaFQEG/KtwoycT16epvuLyyihWQtX4ebnvH+M+rIA+qbgcnHXAos9+Y3zikG55
qOZ5GUD/05vgpx33JPD4QEhRAJznskWX+9NF3uWeIikGn5oEowI3jrshEM197eUDznlolN0XGRXm
1+0FbYjhypIitEuUv9jezivb74g0xKFzFat8wOiCA3LNO5rqq5BKPgmfL79iJg+O3d+In/bsD8xi
V4ldI5yJHebBtcaqcfDmHa73B6HbtesstVQ+MReH5J09Gwwc1ZByzqPTt0tFMXgYG5FkeVA3qbI6
JBvEUe7KDoQliCEP0+wmnyIq9xLndG5mzW/4lnj81PwwE/iabF250B4wojChB1afRCb456A02ZYM
2NeFljaNKSumlXxUBQdPZHafQ623SFi47RpXylf3wI5JrQSEB1k8Tz+tt4SiZCn5aWDIW3V3vZwP
mnuLkkulwnN7dU1TZTfTFxnYuqd2nHaHQuokPwVx1XehmAR+4rleTjKDNOB87PVfPI0PDO5unZlT
3nJ8HQtU3jYbW9cweoIC3DSsO8naoHjlhMQR9SJPACqj1C3Plsb0iJccF8nqt2y3YkKN0mtllwVY
wDlH2OQxJHjNxJlPsfQ59RB2gyMzb6aqDZ0VsRvROOXgqUPeMiK4QBrIVt1Qq49gSRf2fqGBG7La
U0V6WLjopvjaRQwpU2b6q9YazyAca1fobzuXkGMhHmQxWKAyR9BYmv2SYTOVkTxvP/juYrnHqPs7
GP+sehnaJXAcQCxIh1U4OcoXQv1C3/M6AtfSNWvRRSQRgfr/uQkMQlSvPuRfrjUQjy+pgnKmVUBK
SBIshF0KYEt1HvhsoXFcoDSgmnquluQuYJELBw2K9JBjNpNEJu/AE6Zk2JMHVX9pX0aBz/kf+iqH
27rAnXFJ1rQ3pYR/vlqlhjTijV2/a0hAuflOonqoSKq0QkronENqosfH01wam8FcVVhF1M5zYRK/
XgQwRH15cGeElfQV1BVZE2TZF07tf6sjefMSEg98qkjDmxZgglGiHZoSw0k/KsIglD7L0u4ircTg
i7FRMu5zjlmEMz32fK9rT5FY+o24HlrNmb3sZdyaJe5pYMp8U1/DEUHCcQIyPi/5JWKknSvT5YdR
kHS4/f4+0QG5GLLaL/mj9Ox3S5hFAtoJS2YJGemvcQcOlCQX6aci2PXMTetFZq/nMbSds3YELfkv
1CWNt7p969a10wE9q4wEKx5j5tURgfy2pfs8IPsqERqYX+XlkHI9Mc6AXv6L8MFuBFr5vRhnl12Y
22y+IAOZ9XafuesMI43AvX1V34ppm3EmM+IFFFDlkp/+TMX9rRvNRW/oSXWGU7uO2GxTgUYCTCH2
gBdcwCDAyWs9tuNzQgRx8gFBOh99TD76fq2v0qm2x1wpY1ZkbnyCeJvvuazWiySnTwPGoU7RAhqy
a5iCgF1c/1zlRWUcH+5jvKl4kc2pZ7G2yMgIJOXgkwORMk/NwxTXOLN+XMra4/S6IBeRCil3O0Os
dXBLVIWPYhKFOpBfXY352mZJ5TCPuFKuWYwNINFAzLEWuRLjKfsK2Vfmn+oP3t9IQ+bO8J8SUY5t
lsKNO/HrEahS0gM9yXBdayS3gmbt6tm8+ZT1MhcxMY5bWfqb/ON/UQy2fgrEOP7pSAcuq8XzLONy
fKPWtMbPZLsp8xSDpnb2sM7USOViA5jIe68+qLT7qMwjszCsJTir3DSmTNf9BAxN2QuiN1moO8Dc
ZW0MowMNtFiDIBfptpGXYKEKxOKCEYgysMoBYlvBOZ7IjUMJPgYul4wXQCKU3eQo0CREQV0yWdS9
MhzqAfxJD67+i91fAJg8g9w387LWROySrukXaIhOPZ6gewPJHCe98yhw/UcwwMSrLRHW5EQriUc1
qxImBlNOA4lwU+caJpHg1hT2UvpQ/7ZakuCBF2ZwOJQLwDNTd2iXn4EfeKPnjXls/0d87GgAH/8F
3Mn7jAXOdiVmRH8wbH9w7LOramzkcott5hljIpxIpKlDT9KcbrM6kPh0y7NlH74mBkA9Qhl6FDNq
jESInnRG0iya0o7L32O839ZGO9kp8V66INGd/Pp4SOg5+nf4eKOEiDSk7P5f+32VXygztTo0bnNk
tYTt9ROG02HEQlhtkLLZX4OV3psLaBIccPvoKfKSYyFpvgV1tZORsI9jI1/E/DmoVXxBqDp74jvP
wQKMJn2X5CsiFUjt4eWa6l+qt6/SLnPSwQqtzm7I+LNGEh4UNRHufzWVe+QACrN2eD4NZkQ9GQys
05fwdQEpGjH9KP5dlFeBNjH48W2evrsQkNgZSqvWgI5LMiIDVyJ5z66lFQGw27fJCLv/Kv6jneJz
Jw1OjkK/qf0AuhGN2zRpJdHjrAE98lkCF0iCTjQOPwjlqSbDDHut8E7Ld6BvXusooaGHs6yurkFj
Ltg2FpykwB5YCYa2e/Dzm5CRUOr+TRZJ/C+V/LTtlY66fnZJi3IX2sF6Ya8o6NZeSNlNASJhnhjs
gxVbFCAM1brOnVaOGmSFnvthqKJOk5equ52VUFOcrN5DBpdulpwIgSlT3DPBILdXUjILn1Ed/31B
151isusm/A+Qsw0lsxmuOCRDTVDLaTDoaNmt4ICvCzVtV8awmsMCEHwDNzQXY+7AWkRjZMLvMMsb
AgNQKHKXlxEk7ZG2gW+HzN6wWazgT4VwMqEBapFMTW7B/1CJe6Qal81Igq0IbCrIvIdv6vL9U8XJ
OHO8SZao+RycwElQQ5wPrbxzM0UJiE+XdL80vzqY8cyRv+Menhlf1lfSE6PYHHjOfgGMJWXUFtnl
inLwHwesCypoc5qgm3K5jG+17tuSDmD1RhVhyWKru9UxBuxDJ7K0UmS6O9isZXey0nT5Q/kSmmxQ
2rXRHmgwVdv5SeEIx4xVn24qnC10H7dQJyzyP3cUGW8jqcbBAA9lPHwcnqLRgwVpG+HpRjAL3mlZ
P4gUi0ZB/hswAPzK0b+O+nNpzJWMNYm9Tg9DemTrb+vfgJwTO/HGBq9WGmU9HYXBsMm9ZWkIgGSd
VmsyAaeNIHUNZc2/4oMid1J13L4sfINi78Obb7B1/XjSdD8g3aVNRnubxSp6y6JSxDmgkAL9j/eC
rApQrSNe1amV4kDTi7Jf5HwM/3QBA1AxXFbkp1BA33tRnvqzRyNC8Z4MgQTp7uYsqUZu6T75iZcS
VVwyOOBPC2R3ADf2PGlQKPzLTvwbGolllmUMge5IaaC7PBYwWhDN34DHSmTQaFxf6iuM8s0kJ1TC
ARMizY2N4AnLnYjnfI7FWxYOc1vAXPlfUm1xhzQmwvRy14HrZczxpBJmKZDGR+cuv3+7c1rsntjc
NVHPW8UdASQirNSzKmTr9oh6Vc4+AVutiNmh6VoVy9aKOx2Ik/EyaSxvhtvA8tPBP+uDYoy0DL90
BHQptSiYfuxmIH42YFgf4jt4DSF6lhx1ZWZ2TUJd4iOPShCcMX03TP3gH+j+Bp9VfxvqosICZAjz
e4v7PKDwxxVMs2GcvhrAR0rBsliQjq3NX5tWSW6tEtJXZ+cfQl9uKQGd0OCzzFGunpwEzO/PI+a1
KBYndGm7ka15kfwHe42jIdKJLy3dcegnCJOaWxg6Hq6mZpAShKu9/wDVwZ2Os9jhgHlHz017YkrZ
cdgQ8XnB9Xg9p/6A2/BxDWQ1vrSWRQ9yHnfSsrGyB40GuPioGGLgonkoYvfNgODg66lWhymvIWjL
vpDNVrEAP6OMy4zVQndFYdzNdqC4Ep7IRJjYN++LwnhOoMSaklH6/reHiDTuOuB+U38M9DtVfaKC
yI2rzRcnGB4Rn3wnwYJxtWCOL8c/VkiaUc2P98QYkcp1/lxxb8QJ2/SmQ322XWd0yon1ESQqv0zA
nxyIosJRQ5hBFGbotMp8pVq0cKY3LoHz3MYOmNhZKW+PZ9Q1XUKFol9IhmfBFFz/0slaXMJcPgt3
/6AQ7EkARErLTE95mhCdUuH1QRUV0mBRwMUsBY142GtzJVUctFhk3nYYDiLbwhuf+Z1VijbeRtDR
aIiv77Rx7QPZKHoJgIkBubixZlU5n9RgaGgYsomOFtpIIp/o9UiF2H8QjwnuRJwwDyfb98nfcAj1
/3Dqzk1o89Rtdzi0Q9+zLSwcxnE/WZ7U5GkcEUKhDm6ULg74p+/RVcUm6+P8nMDk4KL1HyWw4d26
7iUV2csh364s8bw3WBnSv2MnwGy84N0oSYnbIB89v0b7uY1EyBnKQGAy+JovHsTv9FrXx+4uWwVO
64wKID1T8cj5Kve/uPOrSDMemqsgitdYJIaHjY9zTi9IVUvgXRuc42zFekg+Ka0jo3257tdAPx2E
yYmOwYxe7FIZ1Lx1trFWaifiQQoGFxMyGAlmmDLKKqE6W3nvC1ReRLMyH6ZFBXJcO+n7PwElyuQq
pY3A2iYP7Flb25VhHTCzHua5qO6XnsBMdAgYwfij6NrDjuK7WiFNzLrgHxIq2NwKx4u8BGGsUXPB
9TNmNZngiNYoVTxNzB3pyHgzpbYfwyInu094HA85I+DbhNc7TQ8oifMG0CFloBQeksKztp7h8g2A
mPyyIDF1UP9OU2w8EAfBu/X8TOt1TCh17wYR+fncX6C1CkCdlSu/aoE4ZQDpntyq0c0zB6MYRf6h
Hrn0CF6kVa3oTHdhFm8Ymzrd3at5vqMG/mTSRBWfSG+rExRLxRXg0+VKiHEa7MqRE8tPkRRDjfqn
T0jlrYnmyyeO+2Oe14jkm7jE+G1PrGyqJ+Ej+SRx3QgOhRz1y9XiYfddKHBDvOvwQSqcJC/CMRfm
xGY1xnql9spSz0kjhf7x8+cUf7TVYLbEEFyqlus78k0nXidKvB0QmwZaLCS+r3uzo0nWDPT7WtHi
AOrSRyoPALs+MV42iewQKnsXvlRZIA2oFSDRQigUiHR7+4NbKEtGGSKmU2f1CNGw6OtOQF07ejC1
M/17KG+Mjh1nYYzRwk6Tj66FUZd4Ij68Y0xTvse9hW/ry/aHYfRYFcTElgqm4O4ofGVZ3KVfl7it
Y0UKIdcZ8XOvB1wgkE0aTNqtw1ai0CVVicoaVALfFRfULLPYdArnV/8PQaDV7UgxXV+Kq5EyGFxY
FaWfvLsxM6k8Un2xmh5VTpgGebLkHmNPWO9j8b852xAjDxho+j3hTF9I6ONowHs6R2Kg5qZ7I2b+
pHTpMEKdXIl7sMvM0oLtQIkqgICfhWX/EKADIJEwHEls7wP7W276iK/9G4OnfdeXvHzribRbjEq8
VXYmO0hdIV9i/OqgtrrkN1baC4APXJjJ9NH2S825tq/JV/H/bYZhdaOPgv59nmHRu6gZW1mharI0
IYMnSkZs6BnnrPgc2HkNvBkUlK0LUNYRezzcLPhCrS9wR2BT2uuIjrlD7uFe51/TPI97EKSfqRJp
bEBdLnkYwehqk6txSiIFnqeen1qWmKZL+t3zq3iTVFv18Ze8iL7yqq+ElNg1RqztXV+t3+4D2got
DYGzcTvShuzX+/js07AZrPLfhzvQpqqDZbGgLUSCLXe8vj/LIVSa2avZDOsbzYpHqxxnM/Y2Ffy5
1ZuQ8n887j+pJG1HI6ieXNL3vXWMKOelsYY1nEoMeTgDAdPUQ8a2eqjLdUojZl6m0rQAfiTaILVc
81AafWwzBC6ZHO1H0biRFic+3Q8ABxkAdrVUDsKMFW+DvopWeRizu5yRBOAj4nr/TF9uegCiG/3P
smLfuZ2RSaYDhwIj1GEbvmlt5Enop4xI93ayqwkwGRdp+vhJ4e8qbKpZjNCaurTCbgRmtG9zKHf4
oyf9+qHPhyAoZlUuEOR6HYxNISPG8thMM56GZjZ6E2Akk6lH5SMdD0F758UQ2tRSLDtsY855uBPu
ABUfeE4XusN6yAb4hrcTrfDexHUhVaV2vBW4ztLEdjBZgapUaoIQGK8XWenMYY4rGtYmUgxkUaRO
L+dR9DHJUeQWNOteizmdJJbvtWKp3FVLLFHuNIl5/LJsWI6CastJVyJmCh4bc4nr5uLICZdtjgfO
LVuzZ8bDIsQ4ghFlPWGqatrU2gz4BOCrVoRQJte4cXqZ8TaBJ/PPrmVIrNmTmfvEmyvEj7do5hCg
Wfmo641j36qC7++DN+X0TIIRgvPrHXFwq4RswsffmgkvqqE0WDJ+si902jFNCK4jQmPrUouQl9Zx
e/pfDhToiHxz2hsi65WtFECKmIsXV+4nhg6cOyb8XdClD/s0dRuWXtqGAx4NGqnDWyFKpYSNwKve
+bFY4sltUrXxofDxkcP77B3/VuU7XhAUFUYd/TjHiS3V6MNr5EG4oW9SV+APneLk0bAlrGeqg4KI
WTSNmaWRKkJ8w6siEiRctTBfilTNTBKULc0I2k9xF89wtV6/hYeF90XwFmIHPUizWnhhTNtbBf8C
iPF6v3walTFU+aJWoHWd1vEaq3FMYtb//trJvtLBeSm/CGueEu7zuW83Tv/0vhSWG9DgOGTUQ0Ou
ah2aT6Gt2/i6/rviN6dxodTcBNjFgF/wuFaU6idIzUdDiaI+l8ALPAykN2JKiDDVpjcpzMDdHGji
0AoHGvVqed9XqE9qUpWbh8gLMmHi0H6A4ybBvmwjQCXvGuA5Mzux2AFRrEk3b4ojGqYqo5ngj9MH
NJoFF7T8Q4AZnt2DC2u2ELa0Bt5QbxyFNozoWs9J1OIkVrTfN0GhgilGxGpstbVRDurIWki/Qj4q
OpN0w6iHj/NBZyjx6klr9C9DYJX5RxFr2OpwtpZWPXAn4QHnlK3Y7Epn0hPfc5jE5yymXRrUjJZx
qgsJMigeXXXaQwlH3j1xN4zHn/n9yzwr8T67PqhD3kTlOBiKMPHeR88wuXfOq1lGGxbGCrytnJdb
KSbJT00F6I2g4Mpic8jhgpJB9eAAWFI+prtKXWnV69VogzJ2NozZc3J2GTswpZXVBMYT/SWY82GY
8C6CSBbOixrp0xU7a+iqSjoQaJNwiRvdBSuWfXuSa/47OJykS37UC0vG/WILd/Ym6Judk+tgEGiM
y4olKgdF6W5jXYQaZJC5zvAtHIr8gHtuXhj6W3uM12+Tc/8EVvw0G8WCMrP1FH42vT1ZQIvxqbd2
hMlc/vn7nAx0xfWJmRvrtSmMh1D9YlJItT0ekE9nRyYr7OxQRVql2l7WB/SBEuFTmxv1/rRvJiCs
c5ZKG3NNMeg5NgUe683OhJj3m/fTKIJV7fdc8oBwvzZHK6DvbfTDhZeqPb2/WrMAO4/ypzHKhSmX
dStNEF7f2FrGRbpUTeHx/NvRr5aixFUqyPfytJDeyIQq9s3phrqBnDc5MtWffZIKvGINJFa0oe9D
+QezjSFvqmyf1eG8rdEQSl5WoUrxyO4qmDIAHGBEtn3N9FxFi1J9SSHZRzy+rcVD2YRJCmDroooX
6r66tF3r+U2UBvAsmp3JPzNWzARVHYc3WhcZVSzLfPRiFQe3FCbvoX9MsC6ixpyIcqV7OZACYgBs
Aop4cWJA4gWmW0owBhCZo4wSG+hQKuOv5nWOln8tEUdih1QtnPObEuZt0rJHdKd6am+UzldDVfJv
2zO3tQ9vc5GY+uSjYiDekUFddryVa4T/fQdXSbEO54Zg6GIgQkDmJAbv7NJ8wsg54dCYIcBs/k3Z
AIk6sPpJKFcq+V9NARwgqbGIzrlX62VReQg0OjgyDakerXPWvoLgTV7lmCWvXeRDgTbIW4HXSwgU
0P7NdqUp5IYHZtMog3K+/UrZcdJMRR5TO32YRDppSs+RjNf4Gn36FXQRckLQNXG9eWipxGePoeh5
9v8yKc6CWjrRXRUjiHH6i7YPhstha1rFnCHSVMssow+n4z8JEjExSOaxpi7KmAhGG+8SGILZ/C7v
Eu7t59oEi8PKhmEUk7lodiR1zOQHa/HgStrDKY58uE6RlKQ+1ZQAUE+jfzTU04J9W7LTkXMnjjhT
vZ0NvwC2TvrAufnF9fXd9kFHU7cnTzhh4mUFiHIWIzlLwcPWU4CnBXC+tYjSDVaL+InsNncfAv4Z
XaQO55Vu1ue7qfjdSB+Lc3whb66HaBUzKHqoWmu8zCh6oh0N+oZ+C3brvgjdPnVOYhyFx+4NzuWA
Wjc8uRnPTeriKBB2HmG6DhilXpI/TwnPXYgXjZjRLZLMNNVzLWFMuVX3RNtMQNfK2zmbZ8c553Gi
7ySSaVrNNK5VSkg+SArBZDfbsG3RHgkIRbmt5o7J41wSD1uhKQeZBqG7Km0YYffS4T484BWrPjO6
IIeh+cas9N2+jWVQGL/y3NPIHjIsrYHPBogdp/xrWZew9Y22jXsmbY10utj5xkgb/rlqzBNoBOyR
LpLIgyoV/0AyhItEnxobYWiHyX2B6w2SzxuESzB9Q5DEnO3ePVNEMQ8ONUb/AeMkb6bkUsEf+X/L
QSVjr0xf4BpBVddTlFi93JX8y34naxbzaFtqlaq2XOTXNuZSemXBpxSmc3PxByzLPs4TAPKAmqFI
4M45+HLpcG4dHIFynKvZzNhuqluMeto2qrY1VwYKiuE3N9THQDOmNDvFCtprFfRi6oRNwTkUVC6u
x1/RaweArRGRhwMvaW0tVKPZ3EjfVI+uZqWLaorkzUnynfal3DNPNXEh0MwTGobgwr6Yp/8tgaYb
DEmfdJAl80zUhBEGL3KBW2wU3K9CuSI+phXCZtatr5hVuvW/H7kmCS2riGyaxPTm4hH2o+FhtrDs
d7Ojg9J8uyoAGwlVE9I5XSChlKAADQi/9hQ/HRCSvucUBojC8rUCibNgLvYMs5XNX+wrnHZHUSDf
sGUYO+BWs/N0Ywu3gIM0vebDKFnfTU4HJ4Pk/kjkq6WvGIKFDS3Fv2ldVcvvldGX0jPprAwz//6w
KS/8+kA7G3enAT4x4T6VSmenB3RqJQEYdwcsLWlrTqhIfTfDnGh9M7awKKlCCW1tDvx68S57GaTb
BxQc0w+8NJJ79lBH39WOSqt9nSdpTi5BKC1JXcSc0e7Bfhe1a2co6BSP1GNKA+txAKx+0vkvuCb/
DuZEw7N+eDwVTUHG1kBwk/7CRmT6RjNg4odetBEyUpMtHEovdd7pceklpLsNJCYeKoQbta21X43q
SbIwrpt/us+cw7EL8i9us0FQiZSb0MGOR7m7Eu48C/ZU6qBWRm8sighTvLdwDVO4PXOG0JD4pyXP
pcmlfbO6LEY37k9wourDxB0cornEm6Xvyw2oR3/1SGPDajBRtTS00eejuQYmYn4n7LPICwLFPwdi
LVcMDSZazsTtV6s5Eg83y9lixuBc4md97r6aVM+cxOkXMORqw1XWEVQG7gKpzW2dmHmjXB0QhdJ9
0BMJDw9B0haPME6b41xsdVKagxLs24xxmxoAoTfyuvyiVKAKRmewQgCkwNGxbM0mpe5+LVVYisDr
/Bk9/OaLawbwUfS1TzV85My7kBuGP58oNi2gaYb6FAZarezDdRj7bjHZFD210VV3DW9jC34liy9N
SwTbn+zf7y04FAwwP1v2fDJSNECW0hTRkKcKbYfIz1O4QjMVlA1cJlX94YZeC4Ca3SydN/f/Li2D
0WGyVnl0TS83gPCh+djCvoKyJoeMOnTbJX+tXE903Sr2pzJTKDex0uIMZNYvPSZLlXJW13Cwa8i6
+CikzERmlGGx1i/kD4ZM6o+gyORyeXc+6LxAwGXDcFdLu/EHLKTes+7OUoEgfyOcpV00i3cXzc8O
LQqw5HSJykzRtPdlvCjYPVw9o+XWgwcXoMRKR4Y4wJuSjVAigxi+NDCAkKI6an9DY1HWgCl0MV3W
8V4RrfEXr631MVGKHMc9UiaB8sYvCkEwJLnXqeyCKY8gLF63rUExwwxjXJjK078Z9/Wtg8ACfXAR
PGbrU8JFAgcMPOi8ieOMZxFbWtP1Y0sA0MCXfC4RJWSPPidqQFd18aceyhXvkvXz1b9NrnayMpnS
AVWd1Lagf16ScZwqg6m13ylA6aeoSqPFkHFsU5MbHdRUMv4VsEX4DgFd4TW1+7k7PCaOEjI/5iQ/
/vRfIaukVFUGMsq/UFZnKbRG1V4E78blHNEsqj1vnBAg55veDzt0aIvIXV5TA+wI/GIC4ZgWGkqf
bkqTX/U1/I5ifRqm37QImtuXa8EjINTeK8OQVgUQfVN9W/X70G0y9dyk4DTnO8ZToVfSnH5cS6Ih
Y75gSDlIOE3uPpMVDFKNZCE1POdFkAsybAhZCqSkn4QHGvmPeRYoUh4rJhaLlMqVz64Qc4TacyQO
Bstyhe7pspKR9XrLVRtg1xbA15A3cnN5jTNEtx/wSl56qaOh3+WlcIty2teghEcC9v0XfjOH5ZYr
lfCTCnV25KvePcWikYouJdZ5bK2dxIHSxfNzq6RIbuiIKjmUC5cLBwhluC1Sa/muDdU7xC+SWb69
P6cmBTZxckuBeWA5bhedy17JKBqay2uFDQvcnaa1FhaAPeWw7lBlGJjcbVL8Oepms1FPGROc4g0E
o5WCFQ+al66SbeWYVzMNs5W65nlvOdZJcyPoQw6VrruR6l4VnsL+jMOoD7raq2EhCQpJc6hYNeSV
En70Uq+MsRID+F2c+KW85dIIrQLIBwS6o2sLes9fj0va55xnpE/5Hw1u9U7IgDsYqDMpla5E1cJH
nPJ6Y2YCzQp/2nGdBvAQZUiSdibHdaDzGNyToSa/StiOkIQEQCOEA8D8gagJmKwcwcf0qKr/+nF+
m1+0jZTD3tEcx64fruKYtIwtak+1/BLbePK34fvAatTm9pIXdQNSPJ7PWWYGX04i8XbNUWq/Ts1d
j5NxGMD3nC0Vutb1FRl6ssjk0lqpkFTyPctU9t1UTN/MarwWJWXUbd7Dwa2t+Y8u8RLM/eSmW3El
lzOPIBTNza1wxlsWTjvNp0fgHU+s23Qq1nsaX9UPvO6FYIXf0TFtk8EiqTzgZPe6dlNKbVXtUXJd
3th8tzuNYThhShPFdBlIMBIjMRcaG7cKyORvO0X5BfO0i0s5oiO07Wvt+ebBhJ3CJpbMVGaZFeda
i0Ljj3x2DOrNKFuUMERdXCsq3z3c/X2oPmgajevZJCcJ1lQZmFyJhZC5/y6Ihzs9u2LAAhGsCLt9
leldaEWORd19fhbfS2uc29yRsDTYqy/0VJcyC4ePEH5K1MbC2hVtY/bx7CEcNZ1iXv8nyHAv4L8s
sxUew66ij1FAfo+O/jmvtthS3B7RdfBu3q/AZWwMe9k0gdsrvGikOGaaUDJ9eB0LOa3stVVNZS6a
uXo6dSwclgePElgMy2HwT5katN+w/G/0rNiea7OReHZsY68Y5IWXoYxo81/JBhJB8N+hhZA8PPPS
2j1aPghxBdUMj/sonTFyJE+jzZrPmnQDHxdsx1e2RaTiw+M+Xj2fSvc9Siu93d5zrnH+bhbQT1mH
KFiXfb4MyXn5uTCRAE19lEyZTXcRhPS1eUtcufYIqvsZLZ51psfnMqiO7L0vru4fKG6jkr5nFqH0
tEU2xdVXA0Z2ue2Rx3HR1Cmk12QH2C8HpYvyMhMwmlxevqcmR2BEri51V66cIoLA8EBX1cY0Gjgk
0hc8buaz8kqQD+/f9QI33xHxNo3prKo2ZrEFaHwULqjyEEkgMtNhueH7D5gmU56xh6zHIV7cjYxm
poiyKYPVLa2j1PtbTqbj3zC0Cjh9/BWsUe4Ob3A4UfqDyA423MWiwB9WtbCV18qIIl7h6OIyawCZ
tcwYvW1Uf9D8C++Yp4pJuNr0NEPPl9DBqRz0mkEiXr41TGRLHMkgaVJSoGHDXB7/DtQFn4zQXyfD
JIRsd/c9y3HiQ2iAiMT0Yn3tPq4HJW0uO+q/RLDiuoK6ZGnCjT9ScXy8zSBwFniOr4WiL2pErmF3
HdUi0WTjLv+LsqyAV3H5Kr6eJbX5vNKmgVdQhOX++LuJXn/oKIsKPj0F5fyl4vEALAJRo1NKkPNX
4Jj94MpxPmKgMdrhSHFj29hgmydX/SP7XT5lDkF39pfRiiQlvWSeD7MDSJHTvnENgFbDi6TYAWlL
uYG+36UbqQslBejeBa5AdvNETuQRiItNKSwNoujdqjokuxlO63DQYpcBSpjkuPL/6T9w3YrMRkZo
b0ewwRDChA1BqBV990jrU9vAKv7skUVyJuHdGmcHmznDoV13yNkUChaPVK/+YYGwCOX+Wa5L0pXE
7Bs+l49jYhUNtMBRTst0goiTl7pUvVghmnIIZij7tWLKszmmW9c4Z9yvMkmiMQNua3M/UkH9H78z
eR8q5Mi9UMdtD4dvgLb4np9g5Ki6VepxGB9q89hHSloj9kYVTaI2LdC//xREaazIxIe5pTgjRvtA
lSUGMejwWdW3XxrFcuaHNlOegAVR0DvNKIad2cKWetFuweZaTgsU3D0AiTlmYZvV979dQ6Na+Res
3/T4zvTax5Qm5NiXM6SJuug/qPbzODGrMQ9kTPctmrcNc3CKFwjR6yO+TUr0hWocqe9Qznldk8cv
3CmKjZs/5uvLoHnv1onIJKWMEa1yVCQdFJDUbbjJFKcNx35Yx6knmef8acNs5TKpDuU4kZJgPlwm
J5Lo66ddUhP+oGoN1867hhh2YSiGd7vsAWwdJfi+a49w1laLwVqy7IpDyYLJxOGjaxrJEHT7//5z
Ty9UhYqhyi6Ibkk7CLfs/ooopupj/SuW5xykaoy+06FYlMzCfdpLu0ngf0ITPLKgLIbCB5oU4tX6
1oqzsbezECBWCWYhpfNImGVPx1TjicDbl5RrAScq4nPs9FRITR9+Q0Kl5NM5AKDexq0ZfaNxD2H5
T90QZV2Sempu7E3/48gb7fkjJoNHkc5xKEmSkCbuMRJ7NxRtp5FAutth/yqbSrJZ3/TQpfMnMB52
b8DP7aAEN/9JqneHLj0LQ+EVbvmy8iV1p+c82QcUb6dWkv4LePZYY91j//zUdafWj5KQ3NoNn85u
X203QEYbM3+vW5+fxrQyu9WhOfT57c6Ns1yc0PnicNn2cCJyou0G5prsF7SZVnQrVUPav27SjP3I
9Etsef1kLugF9xn1XThjyxGOJRvFvd3B43Za+fN1w45Spd2nfoybjGP35stKPONza173Fn5QSwKC
DAP7vdney7Uq4GrpO38aFHSbNoq65+RG69fdc6DXeP9KGkpLslh1Re49m7fOuIuSPg3Wcv+arAZv
cVX5X/fN0yVo4eMf7Iyd1LnKevBJVGBs3uNrIn+J8J3yNBiuXA4zEEx/uuXNwNPAmu4HryACiJYZ
PqlBMgtxDmJymu1zCuO1waXo1JYo4BdHuTu7H4MoRNGCndcfiCJTklXdLIDK/BuMBC2I5hDVeDaD
N2Ayre5j1jg8WQ1lHgfyI4pFTUbSBXxhqvCjM5NKroadsbftUb03amoyfjv0rt9tcST/Q5oke8iQ
TpKEQuszXiwgD0NG7A5p1++ALjsHhEbg3CN8bahABN6BhFQz0bfz8Cevhk04Jc53PbbHtR9plVWu
QbHtSbt6nUSNe0RDFfpU0josedUvhbjqrgbKrPJvy2p9fCQjpucSPHsr8739K3hN/AqAW7kICRso
NPLn+NiVTRmOoBu10W4jz8uhv3PxaRtoJYEU2WuTSbWENx1bd3mtF1jYdWMnwJnNnf6/YDdTqwGm
HYRMGPLNLI+JLlyjt3yZ/Pxbr3bnfkNqw/4ld6yD6sAZj811mArJRQ2oT5VVBOC0iCbp3szfLRj0
k/1CTht1Lb6Db8PQ3tgLaH/0Yj7kFBPdtqA5SItVDtoOX+PhVOaoyKkScbF91liEGWjh3YeMM4IR
5gbCB2IF0eilB+Ghb78Rf+JpIEqUgXzTgmHawpxhM6Ap1cqXnCOEK3lAf9ikr2WtbCju3kykRrog
PbF8UZt+aBafS5H80ymvj+rOi0DeLplf5+sXcaS4YZMOXTsWjwCTwjb3q3mom+jHAs8x1CphudXk
Urk9uVDcOlOykOMef0ejtyo6mwifFj7S0aYfnkNppQu3PDSkuHuDCMpljW74A/JxuNel0VI689zH
X43frdPFYwAMpL1hQmQT4WPqKraUf4roRGlc3CnFmp+bSkq6pYLkhtiOtTLui+wePHW6ZgtuyCpw
OH7VFZzt2cBvxdkAci4g/TZGw97GOIitW4WQTr4ZDtnVQonOb6eRbZqzEWgRvG88pJzQ1WQQdWBq
Un98+pMytfbqdL3Gi89afjpTKb8y2dUVdHb0G0p7OlPok23Nj/k24Z2nSUjV8Sh78FAUV5IRNzfF
1SfzLlsUIEchAXciueUSSOH7gSkOiy7VI9DH3Qbw4fBFHT910nCJ30szU5f2cibUyktBrOK78U8o
ub+zC4jqiK0SRtM3j+idVCCUIb+E5N1vNrDBLPB/q0UgkM3SewwmoQdqmtqZbWqaOR0x2l5y3xpC
Cb27AOi6UCzj7hc70oq1kpXQv+C5uncfudRjzq1D4Za7fT6Ej9uV9Y0ddg6PiXz38kta9R+Ja8wj
byM7wIeyusYSS3/TEN3Nx+A5st/YdNw7zwe2Hb5UeXG+D8wvgJN6eOLWVQivspmUDOFuJMb2c+wj
mW0r4xl8ZBbyz4TM9S809JEp7yMuwypbdQM4DDzuDH0cIRl67sH4901l5qfrGDHqUxCcosqVyUpu
X41J19HF3C8Tyqnea/RMQuRl8jCmPxa3x1G1pZMu//wPwRSG64677UKk3dW5nsoeZSUWh+aSU2td
ZVbODDshSlH1eEl6PhtFZ8ZVfEyV8xNJ4vaGf8lw+gp/qAje0J4ZAFujTY7bo/TYPuEFbklrYpKM
x7rMS+nFbjRb2SRrYYM6ZSS0nAo31SAutgUn5qbxkMYa/fvi8CdjU4H7BiDuK3EnXIyt2Vj4Q+Gt
qarCewwCQMBsVZom5IWJooyBqT7rt8N5tJ5toccmV8n5IcXqDeQiZgOFXU5bfiVfiJNAJwLI0r1F
4i1aXr2wHq1mTjZnVryZJQLCQC6sXF+jnsiEFtk529HtHxwc3LDzu8BBpvubzuYejn2grikNlJi/
XMCV3iPzP+jryp6IFHI1iCiBNL/DcdmrZm93xt/yGUQgMiR08MadIWf1vktlU+HbsTgqTWIuEoIL
TxoVvoee+JEHNYz6RZF/ubWyvXtuyegZnncYlk73/h2Iw+gMBARyURSYmrCKN9zbrYRwNeDfHs2A
8eO4Dy9VR5+8hTFDJa2+VaxU2eSn5/6I/ndC8fK0bf0A33t/8sYaaqLuQpbmzGddzB8a0ak8Q2OQ
pFoVy8KRsLwPUfI0WY/9lcy+5BH2e+goYHfpdS/iP2JCizzrBGMI/Ykh1Zo2UO4L4gostQu9for9
RCe86umqmhdC97jAKmjEYlGuR1YBgXeFJUmiMr9Nm4/KLzD/L0sIMbgabWXfEw0M41PpzxiUhrcy
fKaZ7sNzhw8C79g9v+8eVp+G4708beA6ZPKo/+WO2dlLHinQ2xpDXI51/hgvT4w4lheZPXFb7w7e
bjt/pyyNU2dom6NIY69kxkvPyrlQ+WKS/zKiQ808kpXpID9pExN3qAoHyEZLa59Dxn5Z4sBMw3pG
tvlVe455/bCXCLYGtW23Qit/EMvHQ914oXYu9iXUySAVLd15xQnQH/Uy6uGEBlRQztv3IZlZJdRJ
nnnI+mpAG0bPVz1tu5yDfZnb7221sYrASgS49XE2Z4TtFnuP6HCGckr/LFUMPrrwt3I1qvM7e52s
9WpVhr39vrDVXTzQOE9PN8nqxv2LLBLRJAbjcIx9j4+72kS898mX/vAjg15zsgSsrRb8d4QH7rMN
sOZKNFJ1l0Mxpw8VD4FufrtYhPW6tUgYBxSC8nJa/GmLSHjPv47rn8n/M7+ADgxCPvAGUZzJ1hHh
/2Bsu6eMuT/xb014SD2nFzUdYCH7PiN9Mrx6Fql7hK7o8qtdaH/80OXh1AJtUGS9lyJyFDjKpfh2
Ris/hwTOPc6g5tankTqz0JoMaBWPd01WveMHdmThTnbOIcnUujkuRuggu6QeUiCZAubitOatBF8W
KOOCpc9WV5X3PX7DGYIiLmYMbiFpyJtDSkOYkWU/wfmHOjqLyr/SCMOl7YLNpgtnoMV4AorNgQ4l
vSGynFsSlXXcEGex7ZX9CJRtW5CEGA7vhXiv8xDQcnf4ezq1Cdli3Wk7etOjBpM7Br04TbNw4/9f
//VEjM/8zJ2spNNrt6sb4P9GqZrC61IMxocUQTi8pPW3+QRwLIQAcqfHZc8nQNQyx7SnFvk242Sp
KeVYBzEIqFks4cf1inP1dryChgjVGelGsbd7LcwuZkDt+pHER8NLgSa7yZ7Aih2HnxN+wX3IM0Cr
zX/EbqyQxTuXOKmCIj+pMesZ8kVaxIJPS2MadTpdixbl912l13uAD7cmoBq2VDUdv97C/A8kxnYR
XWzDaKH8V3nL2sqxk9mUFitYfm/uoiebQqZo+4aSUUEC3ibDw2/j4xRnZv+2L2PtntT3CRoU4+OL
r4wcL+wlDrnMsIBdjdLBmCFWb/Yf6JyJqYaWtTUdmGgrwVj9QaCPWPusVT+a5zL2pUdZ4Wo01y/Q
Y3KVDSeYvpLYWhbvTX9CqUL1Jk3S39ybynRha2yPnzp+sGCQAyeE1q3/sU1K8PyW449IEHEuoRDY
Vaz+DllmC7u/NPDRgXuKLX2cxDr4gJTyPji8D4ibg4AkeGXEMC1vd9KoBtOGlQCB+WQDMeYbHiuT
LxegKJHaZ/afjObllbRCsWbyqoqLEn0eGPrCr6KyJltoFEjXshlsHzlrWlGGCiU4P3tlq6VQHKc5
Wv3Od1TQjdgmMmGncOGKHEFf+i3QmYyjQbnYRixPuWUBMPrlrnBU8dep1xsRxQNcvynghO7boB6y
Geku3RhKGBaX845QZV10UxQiSQgMPXAXvMjuocKqzOh3fbRalZKvBk0isa/ZUdwodSlzrxiO7njq
XxbD4sAJEtdnRTIz3tXJd9u2ryxoZoIGBgJIP36pUnnHQ37v7tlMSt45+vPGDI7aZSFhBPxkymWz
LAVIuQ2gzKkUUcSmFsnz7eMkUMfnUpnshK5F5IVzpGtUTs9NSD093rXoQ6ozApTLTW/E6HPr3XDO
duw1wZHpRwBPUOBWi04j6G6C7cDE4/Qx1J0GnwaW8a0P9P7XtEGHz7tB/UkCNRQ96r6X98w1oN7I
GE+jyn3n9pwq/+poCxmx45HmDHgq6OZviher8YbbNn816tnQJWv+maANveN5AaYMlsomhm/alzGR
NoTso3P6gyq8ecogKr3NmExo0jCK4/kebmw5niOf1CeKLIbO4rHrxeS1ntRgxkNMxp49kU0ZVdpd
GcpELuqh+LkCg5mWIrdekCsgyCTUKZaXb2+S+Tr9zUB+x8gOO2OHrD/l6yHxW5/t+UxSj4RGMlNa
9O6r3S80Zi0E/NbEl39AedQBREEojN6rdiqoss4qSdSahOAA4M8mRUw2NMeIcFzEFZAMbKVXmZm4
ad2PETjIW480OwuHpYlNrP6vb0s1RUSA5jZnkKwEXUYoJNbmNXlLcc+X9Wy/xkPeJ6Adkg7E4S/M
r74pJzCotrnYk+4/kQbPc0hSM7QdPDdOV2zTCIqfT07fRvvHl5xKJynORYGv+M0Q86iTgKVc+/bU
xUy7EZ7j8JHSNhopbW2X+iplruRSTdvN5b1+6BliS6f7ioh/jULRTh6xmwRusrG6leN8gpur11ks
HG2vIYGkMgyu29kT5Wd3SNHOO4DOomg/9L2On/ES4qq+AXxCqtayCormLDX10ZwGzcB7mxhNbdGo
dycgzJZ6bB+gDA+zKlGhaNXRHhGPbhKJKwFLzOgNFE1zrbKg2vyNdu60YuEyc5xQcVB+xFFcsANx
5WGN1A8+5usD0gK6FvCe0uWw1HG8hEvPY6VDqZZgPtR3N18ZOI8SJRGsYMWgDJMaDEVb0BDT0OT8
c4tx8FKJ/uKjDoS8b4UXkWfGmWJg8yqxr46BXUvpJophsw/G3SqIcPtxgJ92/hlTVqsjA2myyvZ/
HynW0Iim5RL9TD5FWW7e+60FfxrFPwfB/kr176L1pisIxNnxJq5//qNh4pDznlifpvH31Dwqrypn
Gqdd5pSJSQGEk+aaTK0xrnvzDvc14fHoMV8wXLIINvaYTj4TLkF+F8hlL+MsieB+0+Rwr59A4te3
B4ipXlX9/7jGZ1Mokzu545x0+ZfcZyIjvBgXtcskb2JlSRs+SGYXPy5+4sHBbRPPhoXa/IBGeasU
aXYfS3fw/o4Lewn4C3Jfq+Bn0LtNoCOktwGYSc8Y3jrIcnCXCSD/sSRtw91b7rGPujgVZcRAyKps
9mDm4jUVhy9fVMnUtTxu2TqX9TZ/cSlbdfFTxT2ctXcX8qV85JLU1vlbKZ16zFcbrzg9qC01Y9/C
1q8LdUI7ZWF0DMgtoiMEgb42KWTp7xVTb1KBEQlgBkWWIBzAh5cIhhVNqzngw/bj+UhtTKma65WA
Xw+dTUACjvU738cs8GIQDQEGAqbF8YUjeeQstiTB1ZArzc1w5Vnx8Pe8UH+n37p2hwbKaY/V9Lvs
fr5oM5vlYprhgk2LIq7dHNUJbWf5rEQij0fu29SyAVn1Sx2pI0uWSaO92eQXsFLr0XQS1FTXsoQL
ETUbsUmzR50G4u0VhNjhwzxxbIH//Xdnag+DPZ4Clyz52NkwDhQP3zeVeeQkKEeD6BAEx+bqRKOz
paWigDO2K+Z+xN6NyNFb8pnfQcrv+zboPFN4XKkQduqLPpF9EGzD2lcYQ/9wZ8uLL6TSuWuOtOaG
Pk466nqJBvIE/l8yc+lj8h83rHy8MLUKrhgpcMmHRtIxVs7gkJcIn6sZZ4zYKZuRwWe0VkRGuzp0
EUY4Xc5SHDVnZtoV54JqspbaQ9F3kSG6pYf2ItGITKcAAm7A+Qm9RJqNafl8jRKuHsYMHutoRvrz
GfvAAxbw000COlKiI83SQdG5CTybVxd9lr2EPeUWp1B3DYne3cHNCQbBVfulO6y9zOjtZYapKlRw
YKdBb2HHUBNnh1Hh0ZfzKS8TC8C6O3DzRRCs8PACtQljL4usuoAOHdBKDBTownAAdx+PnWFCcXco
mzHIqRoqKlJBKEXBc9NLTYOwMeGLM7yyIB1lDWOHo3YjK+ksz6dAsFMFfv6wDKQeuKscxqJ/HdpT
gC9VpDwcFgjDSPUH0fkvjCqxWRT2TfPHby9lNFG5Bd1gb9HxHbcoCVG0sFIGsJIJSixJL5IRcoBl
BXngxZliGnMWWZ+OpzNX0PqpWCg9nlK1NzjXR/n+34hUROt7ZyjhHVLfKJv5iRq8qs+BvuIENAR8
RQDt7fzSKus4BwrbUtf3DssYTYJCFmr+mAEYE8pwEwJ24OZvJ2IdA7zuWLo+NDu5WY5MQlSXLMsO
V8GdW75vaoNVtlFRagMr7JLxIdX+MYC7TE/f2h3vBXh5lJIiKflLkRNUxIUJtd9sRRo7Kn7RkKsH
S9r/smjYXWp3hGrO0MzNVOQ6OU6Vgo3pDcxtenT5XQr0dXa5ufamlVnpkwK9w+6y0voqJKvYV1Hs
P+kyuGVQpry05R8CSXuP1bsteHoFS0ZNA9j3jjQrKvuWbuzi2NOBkBke0I6ME5QN3WyVyQC4pa4x
dxpEqAjm1BEpaiustsLYd16y8bF3n2XhWH1GGZX52DHBmZ34rs9lZu0kFpU9no5jQmwXV6MOZ4WU
Sn68w0yMYagVFL4i1meOYNCVJ4tuMKGexK8+5/6wGbe0rckvVSzR5dZRMXJk5MD/iMo0nrkSiYVz
lGPTxrzqtvI40tBlTA0Nh4E5gEAnqS5sMukh4fe8izHQ0Su71i/LF6Q8f2KybpRRDF4+LqVJ28lr
yVtG+3YEXMZCb4xKtL+PpaZrrGYWs6x+5Mrv48b3uFvqs+GOFVgvCev5S1ZRJxCP7c7WjjCfcRUM
fpLGAjTYnmuWxBa3ZpO6BvUctfJQss1tQC/PKRD2xSrOjO5EPZ5Al1eOKwFKbPIH3pTnH3dqI3+9
EOzNLzs4mJ+4WIcwlpKtHe1urLXVohi+EuFznHoEzheRIqtYHeUbT+t69G+pYEnp+61GVslUZbKB
iJgX3FiPf2UBJ7iLHwZvhdk7YRuL5iIMbNyyULkrswogFUPxm+tkPvKhM4tGLQQGi1Zy49YuNv5v
AqMhPDP59grCgSvJx6scPNdk5SQZd65mZ7ZfPNC14rGpxBbe6QbYOsnaMaMgoj5ulNPIY+xZMfEY
7p03ZxVo+28P/k1wYtry7OI3L8OrOcNz9wtBdvdVAMbcnCW0ZrqqYIU8UOTIPDJIizvzNPyCMezR
SRThVc1y7bq1VOorngBgkbaX9+h761XxK8XWGEs0zByD9R9deY1ZUN+GSu+Pov5dSUEMZCIkoF+k
Zv0Cdk9eshVbab+XWmVnJ9JZlu0UjZjC3Hx8aLNHQyt9u7wkePF6uxmSnlOsCd6/nyQZECooEBuA
UYzegh8Iy3NIeo6fh8I9uHi5R4gFDcK/4rqHnmyExGrZA8xypv2DApduXrLiOck/Nr8V7mzkv1GA
SoanOzTLpYsnbqH7x2Tg/SbavL87NQkrPM8tqG1X7CX6i7eHodFB5PdPx6RZ50g/hH7loszfFyPt
h2YydrbFs7A+dok/bIG054DUoTgngUaTHue3kNvDna4avJffdy8Scy1hy2NseWujrIhkFwSKDbIR
AHGLm33wlquraxhER5We12SUaPvLrjZpKPJYV5USIjHdrLAOFMnOB8/EdOz582cgN5LpJ+i73/7H
HFcGIJQOhhngMWd14aACcDEZUsoJ+LLxN5otoXLdILNJFlva2zEbnTxud+ag+6pN4O8HLnL8CQH0
fw40VMfoxbO2a5LOXSS6LqRZ2ClqYu5giLtrBuEaj3PPVlMtJx/cIinAgselziujBrQowiGPMUmF
mKD0dvVwQyaZIoLE7K9IHW8MHTaF4nBT2WHsJnK2+6MgvgKVSh1G1UqvP9smKKHy3FUSmRmj+/wc
kB4d/B3K2wEra5zkgD7EFO+IOC4mlobFCiZRcP6tt61Dd4evnh1Fk0EiErBofRdMn+q0MGwC67U3
nT3YBCISEZ11qmIQICtypD8yfD1vUykrBhzkQovGL/O+0NBQpEvyDrrJhWlqmEnTQXL/os/HWFy9
xkzZdKrmA5G5Tv33nNlOzYOKBRhUGXhBB+jpVuE5SMCSKWMAMChVaifIu1bq3IfBrd9wjpCeeNvY
zGJavam8GuENJgXREYWgVx9D0vibhR5eiXYRLEyC3hgsly/2/ELWR0lAYDUdgte2ZHxnTzXh0Tvz
3s6JhKGHfOF9s+zSGfCqslYX5lgYAQgkdPchMgKhZh4iQBH7blIMTdo7r5Trstf2qXCY5Kf+qIe5
O0fFZrO3Da3+Vh5bb25po61MNAt8Fxe+FhLDsatRlGuAu5tmDHDsl6JlubSnZVtaRRMfMphn5v8+
6mh158tPR0LsFOtEHpoMDUTHdAJRUBmksXWqoed0RR+ef94iBV86Z6xkxHI3BbV3hfXbyJzBILoT
9IEGhc/vhRRO9ahdpqrY45q0EKJG97b2pGYZVpUEnbYIGDTxsc8eyBSYtAOoBs9dseg1tAKnOkGR
P3qWtRRertPrmGbwl+oh73QNobiyhWuHC4dVrv6BGPqXOQYTx9JPiei74YUI0HB6WT2SjI4qV1Mx
US8lOgm0q/ARJskSFvce6GNGU+gbE69sEiiH8Ph1DYakdCtH+ivvIO7o7zwnsMxkf/5ThivzWLpl
a66uTi2sGm1hnDxc3VCtrf+3CwuIohMGTDl/WftRiSU0nMwOVD0RYMcgQVBwH3Rb5YrZJ9vB9W1f
5lKYNzDL6Bh8LUeBYbc345RezQ3zX8yem4XgZK30G1G4b6GJGMeX2AEf6CCldOJ7mTHr9kW979t7
fAjp+c9Lq72RaFQtX6SRZARNpRSjODlQML1NRnQdKTptUGIly9mF3UTwvjzmSqj8qAvAXGzS+CPy
wwqh9FThDs9bW3VcaMrMWLa70njj61QdWsRzFyGS0ZSN6HuNoJky4e8AuoD6mJv6fOCDaUM4lqTp
D4kUfApMbBCccRQNg6DubjvVMAkFbeT4r4O6TfR5XqFqrUVIN9KAo5OLPmim8L5K35McTWcjOFGp
0Z8hW7fQRCqKBJRJZxJPnxnsJnYueluKf8cjgGoHDWlD9ztJKWkd2DGTyknvXFX2cqQIZApfI7cv
P9/heO/4ILHDM4q2TVtuhiD4nVaU5Ug9DlqaLmmd3ymkZjuiiANbt1eXZMMyc3GnZkD85jnAhP5Y
3eFOnaSd5DmQyOzC+/HMZLoO82A5ev89RSTdhaRbciicgf4Sr0yW6Coigsri2/TXtybaohGpmT0y
Vf0bf9a0k0igGLr0cZEGm1O7KA27uv0hGFGpL7aflQkM+fHMBRaqZ9+h2flQ+AJNsxSZkpoAu/Rr
GRdskk7SuU9ZekkjcGiVWrCCQyZrIN0PLR0/5rHFzXuntCMNZ5PrvNMnnzQHCnt2B6c2suRE8sn3
UNuapwGgGqCTUwPC0q/jky6Yis/gP9iLJXLplyBousj+RrFU7WgwAdole9yIrtxYcbyBHBj3N9D2
yVgNl0XpaL9ZpZcvHseFfDlVBNSX3P0pajJNOr8i1R9OIAH//abj9crhyecrOwITM7P3USbF6u24
e9OPhx3wZxsg0X3B7FCEeFauBTXgUanPHZSFgOD4+JLddrWjoKB8yXKkjG5qfQam35X/Hjz6e3wD
ws9IykfFMbg/kqiLYh5QHEOq1ipqeT3nEslzduM896CTzkB7sisFvhxugy9pgqLoy+61fa2Eu4pM
M/C2czkk3ZrAhPXGMLP+Dne3W/0rwgOcxUBRDwdPgET4gaD29YORjhkt3AR09q3XB1G+iEYhWGpL
2XOc9vAFD9rRpZ6/39Fq5q4Gul7kFeOTPF+XDtz8W3rM7YYTwvQcdTAUuAJsTbzYH2bJ4kb1vsAz
7Bal4JdmEU80rgzTgz0pxrF23ALI9yHMSzJzs4gAaEjJZERwYIpwmHh1fobZTV31qhYtfgNZYP29
J+iewm20Ix2oWSzBFDQ5lC9KjmJni+CqTcNhH/NQOxJwUFeKYjC9YWTUrUGUv2gcWci2LTawbRV7
/kHOSVMjc2uhyY5olyCIy5tmsFm1p2CsRygCoZSUFwrABT14C2GfxRhfry8oON4D9v2X5OnNFPf3
ZUk0G5U+/vBYdi8FcmyOIySa3XWz9cYenZqVbKcwiWJWWCMeqqsErDQeqpT4y6SgGGqQzhBDNj4t
Emo9QMfnlOoI7H1EphU85PFKRS+kCHHioKuOy0oXI6EuGAOJu78tyRDeU1lo3w3slUCAKs/1tjVk
2w8Ao+8+uOuum1cubYb2Uc2xwDFhcCg1zSvCaeBIQfLW2fpCn4eXF4YPshK7XZmAigE3sE9OvyON
JtpY6Qs1ryUjM+195/PDqB2/BTOg4Xk02CTWmX0dw75qDIHMk9U3IxaeVN56ss9OUXi5Q0NqQxjm
cpGkJUI3PsgmBLDOHmLd0cXWQzo1Zlx8v12p+KD8H+dhDpXwe/5F/+zpTeU9IZgnAsVy7nrbQ7fc
A04NjK+t4L11rB0Fg7K6UN1qvn3L9uKzoaSmvwLLBUfcPlIBRksGsvoEhNpA9+dSX1ijDQ61ekSt
KF+f77a1KLBugFSUmgqwLZw3yqQlZkj1/fwssvK6ZGLS6mAMch+Z6Iq6AqEIJgWbCWy4p/vI3DfD
cTLFfxkPaBPUQDMlk4n7p7y0t6TzjaI7+icUU0r6llsW+5gd1r6CSbAh2fW4smFXwJs6YKXQ3wPv
PFcPGwhW3Au6pgyABDLpp/UmynL2CSWtywmVmCkr6Rg9v1WN4mzP+APXQED68Ksoer4rx9EqDkR5
k5Rkf0Eh3SF7oe49zy9TkvPlWDc5VILsBoyU7V8r21kyrzSgpw4YLC/9/2CAcncE5tMwN0owz3++
+KHYiLm9cMShp96F5KyVGk+79m9j1T6JsE470cewnUfuw/BtR4O4fivrojsqy7Y8zEyRjPmamx42
6P2p7hTblvVJlAtqx0xSZeQriyZciV0cXn1rXuYkM5V6SOIiPJuQRYqck/utO3EopV+/acFD8iLC
9PkTvueoSmvpoE9cP1KgBxt2z5N2L0u3YbVT6nYVqwFVt2HBd2Q5a83K6fOyeH/q+M0m91SDMEnM
2XuD6qoSSZVJ9+qKUibrJkXmjsK3NpZCkGjYG+UE2xzDQ45NNhX64b+zj76k29Nn3qhlzmRUug8+
2OQtMHgIaYcP+SqKPzFcz448xVHQ6qhNZ0dJD+iP1kKB4yjpIWpLAvIH+QeLRGTuzms3i/lWnLmr
7kAL0BXBAScyXwxEJR16QtS7M27fhPvKSIKMq4Agwi1+zwWLq3kvux4El+TBsELVg5jftzEGcSH5
sLutvQssza6VawxYowb8VtfbBkFXJpIWz7VwDXZUCeQvLzl8E+RcGdyqb99XyRYtA4Yj+dAO+4I9
ohKgyUAC91bc+91DsJxj0N2Rr1rHf6olKimaMPPrWUF157bnHBqkefjJcAfOEgDdfAnPINHtLVSL
9qtb6FxlkkPUsvjYdjhrZ5EHB6yVcnOTdYbxqmlPppd4DTYctq22BBAuhojvnxSlFwXpjiYuMHSn
H4VG8UMShh0SfhhO/jrP+Ndpp8hm6sspuDR0Qe3tiDXo45NmdECRu5L8aQ1cxLn6s/pNH9WzaiKu
2UqA6edFDfL0lDdbjjTYhbi89N9kcsYVMXz4CPOUbDjzVlj6s4LJKjgR3XBgNA+Y1QRMss6iWBo6
pCkCTKZ4nU8eTGOvzqhIWRz+tGiXpnMV2WygY4XqcslS6dJm1IDQjyzEkyx1T2z/wpWFN+2BAHAX
qY+nqaYkHYtNnxtNy/hvRWGzGJiZ7Bd91C/O1yN10UUsLHqKAlRQYsHEkKKNMfK341QEuxv8i6Lw
ofvV8b3Q4xT8zEb6wg8kFIQteQhRFB9HaG8nNktMigwXhm6ZWGturUH0AAcDz/oVYCmYzKPgIsQO
cuQEO06DJCB2KghYTkD+d4hlSLfPeXk3zF/+DvxaX1WdDVq5/KWlYJKO0jJPx5bjkXXOzBO5rcXx
PVqS+yNJX3u7GW+Z7MlaktWTT8FDIXJ0QvwuzNqe5WjTbEUHGkCQNn4BqioftDf2MN84s2Jl7nIr
vT3+8TOho/AUBUHaevMaO5jBiZy4QVoPuGJCBUqrfnvvRaQPGwNlWzgW3xNXhFkDKzt5h/XK+UjL
JyS5sgaUAvqXw1HXPfsZgVNd5WpGoIuOecKfTpwuv3QNzJbsuafro2MK3F4yaRVXWtW8w3/c6sgO
ROwsBnbzPEhJz+vFZKh8FRGKsHJ45hYYmUActa5wcEInMyEJoIm+82Y4bPj2WU2u4jtDbL3Nwot5
KGbEEbJ1k4ZqIWQI2ZDETPlIl4Ibdb7o+iNI5/A3MFub/9ZlCpyZ6/RQ3lutXiTOpMgH9wHr9s8i
l53VwkLoI/hJt/pjM/r04CId0zJhGWSX3PFMinDohtSmQUa34HH07/3nJY+RJZBRLvKX5QD6R835
em7HvKKe3EFeyaJP4GpweGd8hco6xymy9c0gCK9OrJp6Idu6/Sq1dP4XbhXUL2YGhNALa4A6Vmfq
mrWalF6zxNG7aawce7Dc128Gwhpru0ORJway1RGplHRds5KdEW8XWwYlQGdmvahROcZUOnEqa+7y
CrNQXSs0wteERwInzzabNMg2TSVamLFXf1d00SobtAy4M7btJ1Jhani8paCiYRLUl3UUhV9j2jvr
wEKi6XW2GrXBLgCAEAXmeLQ/zeiAzu4dYUmqXt7mfimMeA706VPcVDjdKTOyhBbP1SNqPabYili6
BsK/ca381CzYsryINYvbOc4HkiYIM86uDCMr55XPf/Hzbhv6xG6mxqNHSdG2RaX6KrB9pOJ25yJ7
Rd3CKoM/7P6jWASwqh7mWvQNKHge6gHcnVadutKpgnClPCjO8kAznRHbyy9BtjuqV8T+y9LPOC3S
avH9FVmBL15VUPFs1qx8tBnM1FnPeM0VBPsazosjKSmoP0Afj7Duy47/mr0twy1/E0Q3PlLuJDaL
eIIg9Fv+nhrm+MWOa4LRkuCHT6EDF8P9DWs+UUXib51MHINssELDyKigOvmMgFZE+Ed93Gjk6VNj
DMHVOcELXgMDo//dPy/vJAL2Nbgm0yCjk7hMdREl2/HQdcQlmK0dl9BLSglIk5C9hZVaj8YdfvkV
Hm/eufK5ol1qphM0prUKnqirTPdnHDJPcKPN5bIdmZApPZspbBoYqfCtx9W7Cp44U3bZJjoh/YXc
WfGAU8fonjJqzOUt5BlUtrULZx2UJEHgrD1tnnIGsNZ3bBlNh9nI8HSQN/74QyL4YWlxIICTImnz
GpiDZAr97XR43rPKnm/ZzeAXtcU5vo490KQuR4v6bwLNvdWp6GTu+t+XE14yS8VDs7s9dX3gQf2v
EmssCHdQTYsgBHa+Yay7bBJuT/Mm9FWob5JlrEgqi7f11jdhtAPoKoOlFKf4uHKvrKI/akuTSlj2
o9fiEQ5yuHwPp4R3+bZJ743lqswTBhQoXbZ1C1RacfvKscf8wv6orN1S8U8spXaW22sPa8rWYHIo
CB0TtPRMwRRTEePMBmXWEmnEjW5QSUy6w4ITXeXk8zLAEzaFwjGpF+id9htiILYuJg++cI3yRhMh
wGLP9GGfgdSbWfrX08MRkxypxthguJ3MLc/wpcpgC0bv/T+fcec914uidFo9+2cWdedQelk8xBBH
bwJWrTWJnXox5CWLsS+fhLI7aSdxAVKQ8Jn/53HbYexeoWjgLlFe+4IXrSX0I4fWrN3p6aCAAXNa
nZDvUUKvdpSCC6Y3joWLvnI7ImVnq+VFInWTZeZ9ek1nVtFMR6KswaFlUMWSkjbHgTjbXQdLegCo
nu0iERRB6aw47LunqLxBSz/qCdUcIlyzu3K0YscJEY7vkoZ3+TdvunVnyrv+Gwupw2efUjfwAiMk
Bi8nGaVNbbgz9VLhGW0DfKNG/0V01EDyJFeNwFsQDF805Luwh6rU3W+qLAN+bzteTIY/B6S6P/ya
effIp8aJSPHJlUELuKHUBo13rD39NYYUiEMtcbN9lbpIaN1oVqrTvi1YzPs9nFx96PF8O714dyxd
5VVyf1Uaa7iZPTrOvVyPhXkWIUdzvxyYPkUXv26kPpMgNDIcClvButwGZteO82E/rrsSPcRUwddv
RztnS8S1KtbXEIrqPADHjtt+iY6rSa7ab5lcX1EWp1jJAntu+o4HXXltq+uzYsb0pwBkdje6Ouuh
3TqU8bJ8tyT+PP0yAiDnr/v+AYYE2NWm56yzdS1koVjd2FciaEpVBo5mUE72jN3uc+yVlFWfIbBY
GfAVsdnkOVk/o0R1jqQon+Bbq1kRPlStrhGkCOX37XSCkvblm3A1HBwIvhy4TDHEBn+FktymySd6
xGwHJAQNybUh3Zq+lcw89rrvtVYc0CeKuKTt8itBI74xtlFYFVOIyDfFfblnD9aF/GF9GNkldRjI
vzTO7YWukPO2/oM9uuhGjTiAetCf2JGBZfOiOlfmfQxZ/RwbaCp3zAJHBySSrxo2LZaenfHbL+YQ
OevTz9drBYJvzY7itsvqNS5y4Bi27PdnjtkudmFqSWPQH1mQmFChPHgk/CSvsPGn/9gUW/yJKvgc
JijcwJ2MHwP7IA/ghQVUQAVoTrkHAqHV7X33K1VC7VhOvQkxnBb3KoJzFM9YWzoOeEKXmynvey3k
WDPTRM8pvwgiHdt0XXkumRLdjGDizFgS13rPIcIrOkcFEK7LWp+psFfX5yzk2JsZ11uGVRNY2i6d
RI2I5KsIvx3H2pS1+f1/Mep2SZIlwpv/4oQxGLkn9Wps7gG2nxg82wHZFpsQxH6hXfi4oyH78g0d
QAu8MEHN/gJJbR5Td+tw6u4hfCSzi6Fv/q5/c8MfYI1sPHYiLZsfsyW6qWZeiPSNiJ4KymD3Cpe0
t/WpngSAey+SCwZVY/dpdOk4sTUR4Oe+gO6mZP/MN8A/A486L6XjZMDNc+f4KuPzR5uArf5+sDax
kADP+V408u6FVpS+vxCPfMzVtBvWPjRbHOvXR+8B1Gnlo0pxyPNScV8H2g5MKoqf6cUt9h4+rbsD
gwDykuadDeghzgKJEEl8AKCEatkGmx8Uue1cF2EGcqz/bXcl7+GuDFwUn6ODs6RogqBtU6R7qKF2
4aWPKVheRV/YnNY0uxWP4O0qAHhtqlgLi7q41/u9GyqbNdx8CU+3Z3zC6nMuwmsiPoOkJZs/+4oP
8Ml7AJn8rkRIE5kKAuPd0iXrO0euusvWv8lFEBUIXHj+4RaJiz3v6rIwfoCNnKC8q3lJCef+bwyb
oHbQXdzYgFuvUpmxg4ObVy0TeTWp/4H+aHxqgGaJpxPixB5TLyxeThWQlhHkI6mLSZynAv68Uyf/
exBwGHjVJd5DobG7tMZImYMLvGBrsN1J5tPNm6pNkNF+lQ8VVsnrT79WpMLP7ETP//62TMBSvJ//
bXwU5TxuNYCEV7ubB7pw4b6eN2NE09nfMEumjF9hTorEAwQB29pCAIBKtELUMexSd83iwFJ2gZRl
haC3SRVVs8S1mFI2paBNsxTejpH34KdSCldgx5IYgKHIrE2XWafwtXsMP3fkYoOsmZjoj2NJxWpu
vCT0J/mbtx3GxsJbLuUGP+0kYC4sykVywYCcH9U0lGpc14kvOjF6EVpFwU/lamyHJI2NQhigU+aN
ZI6G8mhwsr1wKQTS1GPEKheRv1BGQhIAUgkYXpKeHK8Jj9irEqczUvJzbDDE6najJKQ0qEst1f49
6sKb/Tphp7lYYpXc+dljUytOOo3+ywHUuv95G4nCpHxQwNWRrVni/exlIKUiWdOUmhSQInPT4ZtY
ouEybg8qOVbrj+GaHrGdYZdHkCgt+vw/dUU97t7OiW9C+OlKMKHJQHXl5wWYhlE7xF2CQLYSyo29
FsLiQBpgB2syC1iiYKH7rt13yyhthz5yfZmTimKEYtUBs7pv3StVBfP20cqrV1nQAzuZ9pjcwOFA
3WIGQu/AwUPYaUbNNBpU7LVVNzTOjb5V5oeD+SPEY0QPeEEOnjgZuofsVxFFtkqcFaPig/gQtu8w
6g97a0vHtIoL9tZpBwcYQpxBs7lCCHPc7ZKt8tpeeHdKuienBppUSrLU4wNsgRbHMxf0b2nxerAQ
BBIe3qdi6ZHbbOyJj7lYtZCfLJRGa4VvkbxQfda/hnLNRQ7JJ9mCZyuwO5mwqvfGI1m7Vw/3ipXB
GlC6CdBKZIgd7eI5dO7SSB5lXuRfxY5kWvdQYRypLXF5ENozg7TBrCoxmplFYT3qHAOpR6aK2EiN
x2IcJ4kQgd/F6hcmyDx/O88p3/c2WEM4QdSC6o6u0p4tDtRtugdD9lQ0wxfux1OBXrPiTPAbZcq/
L5PR5C4iQrx7p4wr0L1mLgjc8hFNh2/PaHBFhIfmVoEftmJKWDrlQROLbq8C3X5wC31wZqzvgukB
/ylerAbhTstbifmzXcEZNlASpu5VVLg6sPebrRyBky+UB0yPL1J+nKsSFduqK7i8ghQN/pXFHC5D
ZvAvhsPwx75N+EVrmPHl56hNGYCflP755DXakuHF+FcRZLRPWFUyX6/yTn31iIiQPI6M1Xg4nE0J
P5PGGhEQs0yjB+oQtsbxoeuB6NzD5PtYdNemZ5Myt3hoRY1GMc8IJRldKdpK/C5L3uEpO1+wFPAK
Sj26l2QZryPjf2RV3mw/rpdyN4ZuQYZd5ka3bxlL/ct5A6zXmTkuodfXNgPC6G2H0nXD886LgG0G
MoOVEVlIDXV3aygJ/WcWFmB8b30mSb+JWhokSvm/QHUaL82CB8FzixmuVHQ7DN33warSDzkkYtX/
mgHTtiTZBkw8GHwQD3IpFbaU1tln2EULVlFfeVxqaNn4PHcx3fAooPCpiuo8cYMdNc1smn64yKfP
PbYBwQKgCxxYWWB9TQ5FDhEgvPtotm/PWjD/PDYUI2EPxS7gPtzyak8CsNVTHuIPZB+pvilMduGd
S4ff+LPDCj7XJ1++1A/ET5Z3LIU9u+y4vir8HmXxY4+Q2oiC076cByr3xOQ2hEjaWOXtDbRwkKnU
jwDAW341w4Ik3C6TyCT3RArmLyQcXfA009INDZ6qWPeE8IquKlfBsyRg2D403I//JDT9Wzc6PYch
akRtckZuA6o46C1AtBAzC7uP3J/08KeDk0QJ2Dnq31eXVozwf/T+uNcWsleQEeATTfuuGD8Y/zgN
YOTFmBiea/hfY69tnzDyQ/n+DsyNB1SZNefui0vI+edhh2vNalpd/022FwdXSe72nphyUL9ivSff
0Dk+Sx5qrmUpbdI5WXSZBP6llVDGqPL4dV/stJmvQmWZunCJRzjeiJ9UPv+40hzu0RVsafa9FMxf
9s/87njeddnSJAOqvajHgVpgCCBi5NaKzbQ31K0ePd9twUOQ2vpftp7M7hEkOWvwmgM1qSCv6XSj
ojEh9r9uEigk+C7tNWWJOBgP1icXc82whT17Yng6+XrmFm8KuUehJhtijN9ulNYWwhaEzunhpLga
qhDcDD8Al7GUgCm4v0PKHNU+pBbg4Y/i7MlkTUMzbaZkgYdJknBdN70RjLqooT260fi1s5QOgnbI
MI5OIms+WHuFrbE1uzm7WRn8C5BbEjYDOyH3rrVq3zKhajwFjOC7WqM87e/AmtniVQ8Dd9XcCbwO
h3Rc9rbW2n6zIa9emXw+0uRr+ApmnOU/CeNHeklpq26eU/oorX/m9DoZYFYGdQNeQz1/QD4oL/UB
mHS8McKUtdqLVh/S+CRioRZmrblVI02pngvSFvcNoZ7Y9C0IIHmvHNVHL0bvDOPLq01EN4UbUvOv
o9S0DKHUZEGzwIvQlEWh2iDD6bohzRtiDRA4sqtq+OMZGCC5dpVbiukLo8KzK3p7MBjXooNlsjwE
m2CzzGPQXzU4mEQWIol76utkUbrZxvmFiSQFpI4JT/ZzbCLkVJ3DqkRsMCe8mNybB8Hwwxc8WlFE
/11+1sXArqQ70Uv9PmluMrl7j4U2Yw91T7TuH3NfdaqQzG8rYgis2Aq0SrBQ16B9X93IU2Y2csx+
YntoBrEj0/xSUW5tCSnWd2QHp8ZCzm2axNl4XghHkbVQGZSQgTL34MNA/RMuIzdnmiOJsu7pdCNN
JksGxK38FHxdwUVK+yE+/of/56gI9m2xWwCtJ0OD/Qikib2Guv9dC04EpsTAHulHnFU3vCV1lYzd
mwCKrMTSViM+s9bMuwQs/Iyv4an9Qis6CFdbqZPnVnqVl4mfvarlM8zKnFQLEeZGau1PsP3SN2Qm
eX2Pxr86tjHDPlAMjasQFJwpCIXqrwFa5All/Y6OLwghLHZ22OUWg7IB4jFa33tfHy01cFOgZ1t4
9kVqQ81rIw6C4y0EBv6tkJMGu4OdoaOlnE+55W55oBQhOZUft1HQAJtEDfdee60VGByZImvmVj3i
SFkcMwxHAwtsUoGxjM4xSQee569espOQLFLUVwChGeYUjvTe0yUUE3ySKkuMOf+dAd4yqLw1ZhVN
EfkFe6wIpqWLEF6JC1m/99srih235GI8Bh/38jejtMUUnkalEU+JPBwiy1ZvF/bRQY1wmwzcS7Oh
lIIWXv1DvV+7VUS+Ckp7IRN8TkQftBddip7belzpr2mQveDePDrEEZdTX1bSZWw7dnQgg9jKgrm2
YgKNztr0pnWHwLFl7vBJn+DZXEhT69Bn4Lr/hu90qCOI1ixTFnCeAbUCil6U04HtLpMban8nYzuq
5ZsFZnd8MHHxx05RyiEAQTjBQijIWJ75GPIuY/wHu3KrGc6zf/J3pR1IUd6/vInR7jc6D4vAqSgz
LuCn5ItNUkb7k/eRaR6I8NUuS8rFyS6XsPFPrjwGR1XR3bLyJHsE0RudYabLzxMTsJXelr8CvmYm
ElUcem0vNOn+y6j1IUaK+7dppHS//vaMdjs++7729bFs9XJ346Md4HgKpZzD22HBn33AxY8E7DlX
ItOOLbzkrz8HYp2wCNU7KysN+fqQMZq2OIhOawRUw5jPdne2tEoaOyT5l2oceAXO62pfCY7BIfmY
ZzPqlkg50SzCjw44w/QVqYGnFm/qG7FIbwucJS/Y3ZQhLvxoVogXNGpVYTVvuWe51kCTt15N8ToA
ugdEOhG1mSdCvizBlASbqVJIbrrAiTpbneYmYOenb33qUJf0sq2IZvjGnUG33b24TPn81X5yS6Tn
BEYfid4LVDpGKdIzSIyJUuD+hQ5ZpjMIMl6pYXC3wV2MsRo2Zch9xoDEMTtGSHNFaf+M//iLdtUp
k4elkCtzw64fQqffzvteJSXy+tsIxPbUh7mQKNCXs2GzYDNp0j6k+Za6M4tbZSn8dA7+Gkg3fOh+
ho4+/LLl1eVl4g9Flce1heWCe3RNQATnTHqI9uaRpVTBevKBV5eMjmTsw+NYNdiCRTSmadXAhzgz
MMojgHITi04D3QcPXbwy25YYc/VQhqOJTYMgwLW0tGtZtSEZCrkUectd4R5ef3P9B5hTyLL1sjHw
/MxbL7WiVnbu6bogvoyY/IGoFxOUS409eAvMFCHTf845ZL5H3GLpyrcNLpvm0xnW2Vvuk4U4jdnJ
oKbZQyFNZkTI/3J3zcXXMwb0cOV+dh2f2x0L58LcZNeXZUJuGCaweH/FWILoWOJHlNIGc29pKWAa
7iV9RyiD7gxr1lrl1MC5bb+oWKedI3YZGpVVhaNY9ERthagyPCPP+LQlOmB8OnOl31+ju2rgMFEv
9cPuMJrtDcxDjStD40cjUC0nu0VO32abvGV0NiBv5pCoMvSo45G6KV5gO0hpSaERyY65mhb2ABxx
Dm8cg8HxiLAls/9daTUe1UslD1lSnaFTzMp05ETtX/EnYIKNcndUUBvf03j/1F79Y85uOpOXBcgn
9V7m7Or2Dib5ZioTg/xAge4EpJ+deN0Bfx+cDTwLUdZPe8DEsWfoPHPS3bXXDYoY5Vq9b3u0sW6q
hmsi7zqA5ouuQYGNuBh4Mid3HwRPUfohmZLkJi6sLt8bd/3nZH+y/2SyAg7c+fxz3grRHRGkcr4j
D970R0eahJwwZvfFRYVCgBpJo7pMPvQgIg3N+P574AC5/5QKeQVN/ksZM20jccf/OZG9p1/r7ZFb
OsZz/pGFTMSFcYAPo7BkHk/mKsqlvLtzEJ1ikyYjFWT1xxFEGnX9p2yOTbg7rbhgpFGRTcvVVuaK
ExjalJTG0Sj2jM06kpOOY/M/+n2ZN6Tim8zZN9RjMuI4JJU152vdKS8DZn0EPHtw4Rk9mYhI7cMK
5dnitX6WHddfgA1aj0D6SIPujgdT7HStLbZpUopIHDLbyha96vXU9dbqWtZCvkWfy/53ATHm5r5U
vHk+bkXkthvce0Ojp9HPpVjyS4KY68F784fRKRnICcOqENmykGemTbsbgmmh8YOcbtx1nd+cNOrc
5FG3fovNqfaTupcBSJXKT0snBVGIk4s3vqaIMiiyKX96FpFk1lgMoHYEzS0F/AL6PTNHp+ss1s2p
mmx8l9G8TYtWYKQi6hHzJ57BWwqxPqsq/tAAiL2HIHYvyfFY1w2ZXV2eDvZ+Hww33ioJwn3fpb9w
CraQkOzQmZQkiNhZvCeLJl+9D/QRaNdljmNiAK1dgclkoKphdQxupylKZvzb0Y2hHhw/QINGPcGp
e1y2XqBoS3432ZWrU+Q2AtjX2xpyzODg6M17vZB5RtzakWP8vcIaa6Jb44ZjAT8pwXE9QBoLG14X
UIwrW7QNN5dZCUrjv4fRmyZdOarIKphz6UPJKMQuf2AjfMmjV/bzBYv6u0VkDsnCHd4CvVCWYYAV
AXN3y9HruI6eBL0pPNkqbm9RAxcCaFvUbcJbXNJ4Bxodr3Ur0JdD0AwOKM82kF3QWalY0V/Sab/i
UUkDhPY3u2rVy8dL/NjrheG3mPW58eBhZvybOqrQVwt9qo0fNIor8OcENesU1G5IjqOU/kjwO3Ou
3CXyD8pLB5ownR4A3tZxGvhuK8bT5X4QZIhvOw+m9/F22KLpvQg5de1Wd73GqGyww0GyA/bdGKgn
bJg4mp275wjVJWn9sfrPnKEkx8scG1aUEBK/kty27i3g85J6taGdfDcGlddQZtvjvOUvjlXuWeAV
AL84fiQnmtdC+m0qtxdnph7NsiR0t1WdNsW9Zag1/Jwxe+RYrx3Ky60hkDWqj8F/8rAOa4JAHO+f
V1FKr04lduS8hBxNhy9hlfSwr0g8xExL4vKvJjGheJszy3ZgxKpcMMzBeWa/iU0AmAdvOfKByAJ9
CYBjQHzppZ+JFqaJ/C0b+rgxCDsWqS/3SH2KaLVRUqDijaTCn4qY+ZqHwJYm51+buxo3Cu29UtsQ
9pu5ZOnD0arQp90OneApl/ygwmQzo6/1+QsveWAPYNV7j4bDoI7iyilJuZXKEcj0lRB0c9Pj/wGO
cfIBg7b+mU6IVb3/MHLLxytMI3Rs1P17bbI8L+CLrmFv+uY/VXMwRD6aVguWx2cqyoukxgz03m32
mrcJ7Fk31QWnwAwWComXuNhaa+2Vfvmo7OA/gM/RXRCflnbUHRsDe8xMwpUAKHmJy8VJSPCy/0En
8F43hB1geaTAI78Wd/JoTGolGJxwKzFnF8NW2rok8of3tRNnsLC8kZAIcl1RSy1wdJHFutYg4UYW
Qpx54E97P0vYV26pDxRR9Gf7c8TQp2ryBkkNo3mf0TBGi6NoKNCXvWWC9lgsg5G490r8MRzUp8Lk
79HQl7CVRSs5F5OmNZd1XN2dkcjXShAOWMmEHFlYf25YY2ZVJz6p7ciRB/9a3fbubZUWDXPVknSs
e922KuV26ZVW6V8GFybp9rTcDE+yiZJmTVwckuat6VifNojKxSCgY5v7jkWtLKkJYtlhgLC65yYa
Ikjal0dcOkeOm9lzKf/6ngOmMXLvsbGuYygSZh+hjBsQNGU2cI3/qN7tXLQk8FdLq5L/cGAkD3z/
Wtfu2bXPaNFp1PSjIbzLwQWe/caO+7X/Aw0TzaEi/cLVMZ4GvYvJfW95K7ryF8n/Xd4/Nx8lrEQj
mqg2aCU5bJexAvtVkvJBPSCL67tq7/HnMqwlGfRFkhR/O2ZiLZKZmKOIg0Q9rZEz1hU/pT7PqAOx
0RtsTIb4Rib0i/z6Hn3QFM5BO8PeIMXurpc7/HbQUj8wdku5ldZnQvolqscaY8KunivmEia1P87m
KMDlm6TUxfzQ2si0wA/zjlBiqlFi+egCpIHjh8NF4Cp5CHB93IlVt39/+0LStdld5Zw0CYedcxCI
EUUT7KBQD3GGXKVtZQzD605N85rIfwDmn7vEVNe3Axjf6F72LA26ZmwtbitP8pVRsIe4h/ezm8MN
dEv6UKgnWL/rh9RV20PxWHY3uv7a5pA2OV72GHEY/WRfsoO9g1kosXyPcmWzypcKVQ99DvFidqUc
g19LHTZxqxH9oTQH0s2vLQMZSL9oRK0ggrAKzDCt/dpAN1QSThvNKdfx3iSnlYZktGYFH4O+WEuW
JupLeJmeNeGxN8gOu4r0MD2DVQbdxc0QZt9pP9TqjAL0w7M+YMPoLjUAlsJKyZdRmIWTuw3BUP8O
CkU8XgI9aZSoP2q7owd3tnJrdb0Gx2ELU1Fw4lksj2+YViFetHZ4WFwEPKeuwkSOBsBN6BZ2pBYJ
YHhE6EWJFlkZSO/QehR1DIzLolQwdIUvYJ701dxmj8x8nNeLHhBXZvH9DjgnxawkxMkXY1AbH45v
RsBlKpw1gYU76RdifaxWOb5HRCM3iSCwR+Pr3quWbxjRJX5JVMlSC2VyNQOSizLayz1YypwFy4qP
A9ZAfq7LnvgYLtBV018F/twm9b1EV6phGI44BSNmeHUlSmMTgqF+fkk7zN24ztRAERxWPQqBep6H
gql0AQklauzAq14aM4vZ0ebTLZoB68J0mTzlDEujrSPbrSiViiws7ViEwBGVUWlH+UjrpaqcexsP
tfV7eyJVkDixI/gIfc2KAmnq0MR0Ftfed5rSc8RgjVsticHmbRdygPTp8TGj1D8F9INrrzZ99OMh
E8t+f+4yOCDB5xXAO35gQchk9Adsd0mOUTAVlQw5jF/uPqKl/li0ERM4RiJqY22jsrybWyNWw37/
jBrNn7B7y8emTrNn3kJm4O7ysHrES1gXasWhEedFC1WQk6RfQo9Er/edY99RyVkX/HQACE2W7hY9
2OaMD8lqFnfZySgRT+jmsdZDit3XduXVNhLs687qEHxgELTJmkPEOuScXIVDF9p96xwTG39LHZBt
y8w/xjCa1h1nzyMAB4Z/byJsdrMf7kSBzUPVub9RUlxu3wOLOlyDCNy3zDUXTufka0UT0aX0QsG2
8Rnwlk8SyVujhY1ENuo82GMXAdOLrQ/8RoVTYZ36Mp53TBLHIdgv/r7iVpOTzL+8+eLxKQO1YfZY
zounuWwwkKPHzWUqXAknsWiNQ04YhrC1/wQNDk4sDpJFnTJBVAItykWj5LHWaJKrBZwnJHsw5rR2
QxWQPQCMk9sJrS+CIaDuh3s9eWkhjQZR12x+mYqfFxFfySGgG8lLiZl0flncllzB34U6CIes9qH2
JLh3rzwuvwAhtgAC1MUQaq6IbH0OHUqy6hhP0VUu3UePjwl681ly7FgVDy3LVg4ZFMhAL+wWnfdt
iU8X+nAnr5cSVgqK4vgbqMP7/ZcYIglaMiSfGsCHOq+05yQpxG0pPo0r5U1GqCSoeiuSUcDp2vEH
3HwJO0VA5mYcf1Y7kbluzJNpYDffAMkhqwLMv7CSKTFDsdwRXriGPgpgq9AayHOybXuFLSmSGypf
hf0a/G3LZ3uo/dCjW80MNAHQxXUeibwVd/G8Um3SBWmg2SsNrafYEd+qlZ7QhrN8mc1eGswxHWFZ
hfniKUdH9qG4qZOcguOXO6AIEmYocnMmJXbyUclqQS4l9cMi/37rfYPM9cGDv63hPkBRBWdynrx8
SHgocah26ZUjH8YpWtZ69HlZAWOONjO9F97eRUl7l3mnFaD61cV9DaOfejdbln+Y9rUNQTEwbK83
N4Z/+B0VoBnuwbYiI2u9Pa4x1kkQQgK7Z3iII4wjoUrMslo4Xb06SMFLlVNVzMuLHXnIypPA6UWs
/q7uq8zR6YF4oaAzlHJ4+dfnXAn0upzhOft2HMASWO1jRINn7nt5V7E+0aV9mXVeWJOLo/dSj/qk
inYVGARJ/KE0O6USihRGfu12Vd+23fA4S3k1WWC9yt6CxXY5vSD2S3y3nZo/0q/rRRU/O7lLHBO4
Vdz56GegE5gOs4KM716XcgZm1sUGkKv8u9pLv6ESyiyjKV/KLA4kVzzcTFH8jwrpjquLshIzLPNq
49S0yQgYvKZ/qU/Tmsw9PF+Z9hh7VL5iqR33TpLltDbgSc7ikQebbiqpq5+k28/cm+p95Rs6ChSd
nyewaBOo3EUSkHUJFrKyI3iBzjaITPDSvWMErcJYNLjqoF+ctCQCHbTsxsi0nAtSp+xcB0QwqItE
pjtaMO9udLCRWHwOy6NsYxzOcIP72JWd9l9HjPBmd5M77IuXT3jA8Iiges6MTU3w3nYPTAzyggox
V3J4AnuNy0e98smUq/ack1yYi7TFAxz8OOxQFokyaq+lQ7kBIQxbWNKJdaS28+iPlyI/x/pAOg1c
fro1AyjEEoes2m9JJNHzovcfgyHY0IZb7KkXh8Csll69378QFiapY877uxrwcs89rFRHyAICpses
c+w0IDPqDRLMXaOAU6WkC2zb/CYzcsujQeJgePDNLBn8rZ0Go0NnuObUqKBP4Sqbg7xDWt39M+8x
5IOiBWu08LWyTbsklnwgYxn0G/pOogO1Bj0qTsPhu3xR/GscXkQloQhlCnbi5eLYZ0dv4RfjQyug
eV0/CELTb/fqRh/YWQE85PF7e1PIYBFxroZTMcMIthEnPSzbgRGre9dkm0kddEcsKaPwlcuHXMsS
ExrXmTSYeWjaS0pqal5c/GWlQSlArqWfufI9/b2Kb/UlW7OER/sBFqyVNCQjDmCjQ25njma1AJQ+
gUZM3koTb7x9Kr0hndzWrpAY2OGuYExRCiH/Ivn2RncO/FdADbBiU0uA0eaKTQhiIGgOKjtGZ9ST
aQcK+DqJvaU2/9U5nwL3qi4PBRmAE01U5e5mowL8M7hDbpMK8TABo2YgaVP8zy+Us/wOnTPDY1C6
0rBfnkCcxuNOQKNXRM2yuOPA8OyW17WVJw7eTyyQ9UJKqGcQ1Qe0BPgHO9iSm3FWKUDLsFDfT+zx
T6vInuoE03vhpD6KvFJCaz6p92BYY/UtzcrngyISSlg0F2S2q0FmNIdEYM6CHPWBiLWdsAmLDNEL
e02CqwPd+EDPQz8oa6u/i4WDqWhoUT4CiLkaNKQpiaZEl4O4EWGwGm+6pshyAon3OXsIuzIcMaoF
vrNc6BInVOn2jaqwR6tS8jSzagiiRMiSxGJ4a+BpB1WvCFl5FAitJPAkbgaDRkMQdqE5IHfOId3o
0u3aD1caCjbNUCYj8KL4L4yjo3tqqaS2Qex7aw5LpoCskNLzEqyPrlWyOv31kQL6ADyim9O/yxTe
CI/esvfZ9G/glnmnD3/iBG4IHa7Li5eHFm8q2CH5+hxm0xz+FACL4jcnkFbkINIphXkX/BNhKud2
NswnxR775EloniYnmRTAKoMPKy4MeP/TRUCR58eS94VOtK5hInGbaL7CbYZwtY0bAZmOko3dU66I
cNYKq4k3sP24srNjKTdlPDgWacepZbxQECAqq5DKeAjIfxNFt7yBlAk6K/DMumxWjnADJGKzMqkE
jHcMsdyyd7obA+cmAu/nQlgpiSp7pFziQCiP8G5mpdZKkcEt+uF3Gs9xRQpzt52iYQ1AOffK1RoH
8oiUNdnkgPU911/gGu9BykEMkNAxejg9JVRZw896eNJyCXTEF8KKuDNc4vViLsZWoHTR63VNhTNy
A4PfdPPBr1X+JhGCeNa42oku8qvYTQF7yHnrmi+JH7MzyUwkTYxkv04JB5BpC+bzdiT920bbOPmT
UzD1RBCnwitvr9zYHRZQkn6kUp5KjrycDp8UH4SuU33K7kFloc5YYsNy99yB74e3Tmy3c6Hgfb18
Q+x3bjiqz0PbbUiPHQ7ZxJHt1URhuxINnGLvKspA/CgO5a2uU884Mzo3teFNx4V4rC8PSO+IU0IU
OIEkAcfI4QgVCzzXQh+2DbGbA3Rw+mNprYsVgtmNxm/xsjPZjjidiwz3621C5P72fh+DUG4ymF7G
ekipGQcmZYqq/dHFvc+9sN5WhVnkdVAKHF8YUcvINvGZYpV4Xs+66aitLWHSGO+bezc+pm1XvgLM
lf0H3CLzklTVTRCgXxhK1oY2rFU5+dj+Pi+AEbs975TOr7NAcnsG6HXRgxWHIwpeRWRCOBnzmi2U
EmJO/ySNAbqyYhbhLCnGpQ9FjovWZ1WaNGEzxyH3ZS9AlShF/Xr8VkgosadgrvE89R0qfO40HG0/
wP4A7i06pp06pYMk3cndsdaMjczhfIZEordJmmaxQVPcH5dA7uAqo6EyDTS1rQJ4LXgnQNcSxy/q
cGP3gL0Zo1EYgs4tL5Fqdg+goS+qpGQR+LCXZWTr96k9MmDy/XyhF6sAXuKE2hdrMj4zwc3HA+GS
qqe7j6nVEDNbxZO37h0Rg+a4oelz0f9sv1V2jhaXUg2Ubaww+Hfxcb/qNrRAPs9nb/vPUWA/Rlvh
+RL6PEH7BzF7BsLT4jy11KnLTO7QLxB2noty1QbC0gTZWfSV4SeuzdiIgAHMrb3/4nx919GLLYXH
3ul5Ln0KO18KUq65VzYHg+SqHmgiK7pjudpQvr9B0KGsxAqMSMF3XQL4/ZaS67AGdarIrelOtyZp
PkV2KiWt7BKhwu4ITiBjIBxHHcfMIy0usHOrAk1u5LttKTLFewrDazLpD9TE8POewVPkqg4Bl5f4
VN+b3R/WoL2r6djX0a1z11wQs4SIf9QpQjWuIZxSM5suZzdmlTo1n75NyLf1D5aS2Eq6wpeQgTDz
lwVDr+3jGMr3JMA99LqTPR2lybwIE7Dda4H8DFoMB5T5iumFoMilE8HO8omCqYkuouwUVFCQ5BsE
V9oXFaq0DS+lqTqBGaFM6S/GxJDiXSvg8GDSdCY85TVq36hzr6aXRuR0LxZFhRo1io+BaoV9odq8
pwyEXRZqLLfsEsaf8yorAD6K/Gulb42zTSn3z7yDUgPCKehhxhySvEkY4lMDlp2qDHSqFGcGAPYX
6iUHmUFQOsdwt/S6iopwih+mZK/h+b2ab66SlBcD1TFf/cKuLTq/mtC2v1Hh0t7Qf49NtlvaFEB0
j6wzENlz42fKI97uNDDNW5m+eeDzr884ncg7CPfSt3lDYMs2Sb6MCryQUlBq2Klh5ah5rSFlnkaO
gCe1+DrraESe6ZdCUk2sLhO9/wAPvWZBaP2nKwYwx3+u/CvHfdp/gDo29UktLQii7XPjVut4tnmt
P8dpZMa1W/gYktrqQSk2EUEALqtx5y3Z2aM605lJ2qlfB8lsRLVXl/+AGsaRmxss3XJW7zbXZd12
0cPOyrznmT+1hHEs3jI+sLmXej9Ledkyz5VTcDvrYonGZLFp2iBL99gR23mXj6AHbqGqmSRQ4aja
q6Ckgwwr9cKD0HMb1ExL7gU7VDcQ/vW6q/CYfT4JQiCFr9fw5bnNS6YCGu3FUfr7xyNduhhiNWCW
VSIPr/dleq01Okyk1YthS7b5OvkrO8Xk/JpGhROfOE6saxb2XyOXwwmI9pGAnVi9gohG6i/0h+/M
qh2GN1XI71cVmTZbsIQf+Y9oXfLhrKKO6DJXkAQdSxilT8cHts2DbOPmz/UDm7gWvhH4wkrcIJpo
JhFms2MbjgTFnXM+/DsmuO2LGd3tR8HbWT/cufVsdeAbFQMK03KuIfRJ3T7SCnRsQaw34Z7brCmv
vxNmzg5icaixdPGxjLUhlOr1OYTu8eiTm5F1GmHryIe7mKf7lRcVbZyqTO+XhweLlIr81cBNIotx
nj28d8P3PsNA6UQfzEqEs/LPxHsgQ2eObATUk5bYZe88nnkPIuUUaT4qK2BWJAgRsJtUYxNmcp94
rDZOpvLo//gR2a46m0K0Un+V4mJ9bjQ2wrsjM2K0Ba3C/7t9JCuo37yjYj9chqHm/QSKwTxsWpy5
vr6cV050AQi+hzaWdJIXn0Tf1Ks4mHaLzOKNwVECNHiizi32xfobl6bGpNookX/BI1YCyJzDZxDv
W5p2kUdEPllWHNrdMSQ/BIhe8l/wUORtfaM7+Hm6ifuy38K9JkYT2dcSC7vf9endxP8uf0FXBP0j
+XN89JRy8tMIx1K/ImFlrGtaSLp7xuhNtO6t28X/WbL0mXYdLLH9zTN/UmjgvgmIdv41ji3W3Kk+
USh8qgCZlt3fPAFJ8h1dvfMuE2+vpOVIOd5bueURohM2TdZJAhJXKwd9U4vsEvv8OUMIJNGGZNQa
yNu/WngBg2pdsowacZuLl2Mlj4Y4r5fL4nhgNoTbS3gZICOz4QNfQbl2wtemnQMY2HMqitLNWp/Q
1VOCJS5hM+fbCS+t5Wy8DNLjXOh9UrUMzgfaTB3eacn8WiTIXvdl16Szwky95oVC0iAKv9qp4Bcj
fUCFP8+NBBWiOvQ2xohOERCnszfPjwbkBPCfOallsQkJF3e3p25N02j6SZwKFb1YUb35W/vqsfXu
uR5lFa2Z4ZKZ4V3ozTW7YSoqCET2SW0b5Shd8b7F7y9EqnOLYVRqPqo1UsUyM11mE7RV9liFYnwK
xJmaTTLma9ukhfIE/oRb6x2FW+fuo9t+B/3LU/COCzfiOf5Kw5MxA6nGL1dwHe087OVzeNFgGrM2
gQMlWhMrEkfIMA2EiVLcJ2VlbSDbO95dMdWBOtHaK2C9+/UxZEJZYFdoAJAnH7gWDjxcabwP7a7i
MPHrG2lyS2eY+fAufyiHG+1yU+Ix9qYlhY6yzslzuP8ETeEYfyOcrr/Wosi3aniSsMbGlB3F5HS+
JPCeXf7QTIGVVh8oi3WemZae09o4BVmrR7k6ZKUySGbk5Mu/M+934tkZXDH1Ze0d82DaruIHNceg
7EgBj84v9plEdYNsbSoZwy6f3h5IWJoCl7QHL7M/NuYdxZMRc/HCc3pvYmo1pQvFHg+wZy2F60jC
/m8gc0hYPMXJjyEkSNx/l7xwqhtvzY1wyeVUE2wTgo9Vr6fP0aE+sHnc3Dcg1k5HdOKLUmfCynZj
i4i58tazyYY5Fo9uwW7Lkg7N4Fw74C9+tCWNcVmA8OXxxmLXjrxvMIF9egcugFwPTiXH+OlSccFd
bpCtnMX5tR2wLk/HRogQTewD8P4wD5iI8qZfz7V9HfFN6LPbRCVJtiiykQGrBTTaC59jc82O2g1M
4a37gwUJgQgiqBppYnQ0Zrg2bm/sgvx9SdrTt2s8njOBhhlKN4Z8x6jBLbmwFexBzuTW7lVdJKiB
qJ9cdppXviAudLtTHv1Q7JpeP/ORRB3Cl3qqbi6vYMQbrP3v4hmp0GTqctXsTl179kpf6RvV7RyA
MgzKyZ0Fy4l0RE1VAwk5KKWv569FobAqK7s2++l1RilHhUoj0Qk9MrHgdQU+lnpRyHVySv5+dY0g
fqXy/SioGWcGzT4KrHSAQN3O5itA5uIXP9iWlMGNcmh9sINRCYI+yHSL0z7hts0jmOy5Y2YTx6Q2
XthHkCN7T++OCJtlEGx6/sM3536Lq8TXsw+gOLfLsshEsm0LSK3nZ7Aq3AhoaNIJ/mhUYnfd+dqW
VLUYRkHQk16Po0/MMp5qz8hqbnDSxUctHUO1IMCRss061XHVIaC9M1GjUzq+Fs8j07Pj/Q+Dzoot
4fx/iofDdI/ZonMUEF7Vpc7EjU+sA5DZMgGs1T95INpsq7js169hjh/GbJvPAQuzZlE3seIoqg0c
Wtp7+A3k8ljk2Nysdr2+G6WM7Wd2mZFAOGZSLe0dpMcZ2vaAi3otysSci9EZcAsR5bR7yPecvvOX
YWkBYhbMx9eTdF6ogqmDjV+coqOGWKrHMgDEz04OqrK7E1EWg/SGQwITYb/ciOJK2sU1l2IgOaD1
gLAqc3KcNVnQk8zwpYaiJ/Bdp0V6eqbTl1CgbAXir4F4Gx8z/t0FWrpJEtOzS/DnXpqXjuJiZ7KI
E3slEZaMdv7GwwgpXfvruG0+ciUogwGXPZb3MQAmz62/R1d+yFnKeoB6oarDHevynpdsRi7Iigj3
Q1hsCQ+Uh7ehPoXkQunPryU/UNHu6tDOYNT3P/wzbTo3pd16JDIDWyuzrqEZAD0bYJOD9BGYbxqN
yFNaWQRaviP8H148sxzmxCC5pvJeGi/gRLALlYqRRc5H6gUYAeKsxva6H6aePmsPhuKT4gPIPJ+J
YO6FIaGeXuyTFzSs8gIIRF83I/lFLGKbkTtnlpJI9c2uwGETDXPgjW5pxB09pPLO3po9OCIgERqD
vghvP29380efDQNL1+9uETbBUqZMFKZNOWt+2Pcx0v2U4//btCcxInVw0HmzGcd6hsSfGdBQrD8z
Z3F1TEodnavi50mUULaLtjra7xhIFWr2P+bX640qF1TumegaME0acFH4iX8BY4Rb5ziMWkOYy/8P
iXDdS5ncNhr3OxA/7OxgeJDti/VByz1WUtc0sk5pJPKrDuNkGk/ykyCALC6fml71m2NHgKFBkBVP
CMBMcIYYHNRj8QkAsV6oHYovT7tiufj750rsOZZY1/afxx/kuXmksuUfr8oyELb5wHTEdXAGbqLp
u3gKZZbxJMAoLWB+nynlKZITxUDy/QAyIxbFuAa3RFtjlLwqOtxlAVhbm+SX0oPmSnt7g9eXV3xF
0kvXqyiAsblZujGdSEjOyX+e74NLFrsnIpffzoh4nMB7WAQxHKvXsrZ/Aboito6TYqLXxOnhil+G
CeSWBEbHL+xSC/u9mq3vF3HI+YmXAnE8uoA2fhdscMDlqIUkyzScGs9O3qWzWSoWKwjqaXII47KY
zBwyFLJACr0unOPw4tFHt8WaWS7Gaf60RcScKKK3uQbPb2VotThF/YYY3DXVE9nlz1luJuBSNDGp
S1BZNHxdV1nsnVxvjNppgstIyHsabbRLW0s4Jvu07YzXXrazXmfWiNbRsk/kUrMUAKkoGV3K5NOc
3qG+FtoT8n6pcPPYQ7ew1Aa5kKe7+b8p3Hj/AP5WwPTLnqDZWITvxfBgN17Utdll75j3iktUTIWN
7yKVRz8SmRJPkgQnBg2MYK4s29oouHoRz1tmUaXoLiglhm1qACWALJLaWZ5xNDxNTnxO7iPoo5Ed
ynRjf4nwSizrLHqFRaKLNx78OMmFOu1xLuRTIEJPtqkCS+RTv891y+P7g0cg4RzV4f8ezjdrs2iO
Jgbbv+fWMH6x/m/jXC24Yr66wKktSt8kCjvusg834zXLxHfSiwnVKTVT3hFCTYRmPTmFXH8/SUUa
OScy9DlFt9DdIiOrPgc9c4u0BIrEso291OrG2VC9ncc0Qf28f5iKAMqpeZVLyUKkBMRFynrZmmJq
Rzhm+eZHxilo+LEqYSdQsEGuJwxDDhOsWQ7R9N+t6SU0/HR5DR23kkN8iB0zOG4hRZj7QTj830X+
V3U4RMWYcO4l0f/xjhn7HVHc8wD+JzeqHyr6OrTbhI8/jwdkPWDnDTrahEM7k2ifcSJ4zONKtKM+
HI+t4xtcsLCu1jeSkWRHnco2LvFwzgGNg/5AVh4Mv0iJnzoYQicd/c27aJpcreb/QTF8oqqd0OwL
9EIws+EbUiytkkCB/azYJurs56cxBZE1ZREBbwvRqc1QeI09hBf1VMvfe4l/OFQ+tpdo6W3qKeIG
7dLW9LDDS68v9soNoTsPUwMpt3RNQgRvVUnNbjNQkWRKoJ3wQle/RpU+XQehcz0dfG+2o4c9u+ov
xRiGzI6832I7SoTljPkkv4wwbyuzw5Aebls1qTnu6acAeekTE1G6cTs2JSf2fereKbAQzUqWm+xu
QfLxUkW9S7V3i0gjSpLMS8ceteYGk4eQwBDfVIpMKQgTBL3E9TX4fo0pyplarx+UFwwU+iSLJUHq
ZvMRQ+rab9cVzhgaodRuf0+nzyv+V5X8NfcfyBuCEw88OrU4a1V0CNDSYURAcQRAKEfgY3kZ5HtI
UhzK2YT8/VQi/s2T5svGynQFEHbNn7RWbuzINrdIgDvGc/mNH5D+WQNRfi+QctLP2a/pE4b2cnH6
SJ+gCReiJWRb65SbHPT6y0yaMs2FVe78f8NXIG4Tz8V8hpKorelh5ywHZ6Gp9F3CR3NDM+FVnt6O
GcoN787tmM8L2AhcxD2UeQMDHz71IXTIIZoFJ4jbmRuTSracUJb9ezcuF3TZqKKt2JQ15qkjVwbY
YeAiQgVmh8G69ojzcZQ2tY5wOUVm8TDitRbpTToEnMWbNzDa9eavexD5Dz/GsC5r/cISxnbSavJO
7fVtco4l3P4FE2a/YwtMzfYnQIpcOjdG3h8Vc89V7lozqNSyUy+zcgRhWpNYNh0le61gGcxkr6T2
WElvc/FDpbA3dHUF9az/mp/zy3l1HmdVrjypC6l2LPc+WuvVlJpb13jo8P26eBPMSL7tI37jUxSu
R2KDY+ga6OUjZDEgEadl27mryAOsnXkrvuJY36c100J1CKUqoI24k06R7Wys3rZAuWZhZNjdsLCs
+No+21nm2wQx6yCR9ETuscEsr21F8TZ5I0dYqnq2mJMfajA9rVoVQCmm2IYLjbvrit4DcEZJs74q
e546vZGCTVaj5lZGfrBsjqMc64wPal5UzUaONxg3LuqnAlRh9IBt57bUN6tGEhs8hkKF+iexRtCm
6xzqDtT93YYKg54Jwaek6THjnR07uq5HZIBpvUgsPORInJXLk2mDFg23iw2GBqkOlouDDmtwzdC9
1YfNhN8Y44bNCofIU7VdLbuNLTSzZ/qcn3ee9SkXAGlcUtqaIzPj6nFn9AEVns9ntymwa131qeDQ
395r8UBtto/nZNqPKUVboscg5PWg3xM0pm5yvsiBACZKgHRAc8vH6RZ46seGJXANaKq6cgCYxXqJ
icPCyQZY9LhhC7ACiIm7eAhymKNzNR8sJK1sTRh/R+62ow3M2HsIS5jBhqix9IzmzTnCVCXFoM9H
Tb3pgEht4fNu7Zg4zGkpBCuBHuyvtJkTM9adjTsc4nmxoxCBkQC5a+8R3hPo1CIOu9Zzr0Wc+vaA
zew2W2mMdnT1e0HwvBayUcfc+/R4avDd5exwl11aWdiXQZGYD4Winerhgi46hCpvd+dxNRn9umaX
eHAc+lgTyvn4uk2i58yB2EgegpYQ/SrDAFl4ykQ+XMqO/9oO/6IAANe1qyayYLU8HYTRIcDe7R/r
TiE8X8VLB6HRrSAzkNR4SFs6uDSRmdRvsELHbaw+0ik1O1JmgF1Nic0yYTAaOU7BZtL+Oyqtzodc
w8P8YHEdwHv1v7sC3RvnwZkS6nGfQjxXbBN2yg9b+U5Q3+fCl23gVucXJByXw6x7pfWN55oLuqvj
ycWzj5OyDjtpiKos/Mzd2TtRs1byurnPEHGD8iiiRsS6Spi9hdA+vh0LckmDdzkJg0rBaT8Q4r/g
/zA+kA+OGBpNocWrjvbckr+cFTfIYX5t+D43zzQaFOEUXgSJLoH13TzQIvch9cb7+cuTU9m20rwT
6LNMLpvFCoicDetG2DhFh6/QGIU3PouZq6RN1hRukJriJZ31t0wJqP7mLQV0uMXFmw1qywvNSc34
21o3s62hTa4UUuTEakTh8rcoaJ/EOTaybp86LGGyTFcnPUxVHQXLPpcxx9+SEmFjViZB3Gvu5ZKN
2heH738RKILaQV1I1+JzHJHjNtLxvci0ZjrMmc4XQmXpoVBTbVE3cm8qHv7BbDohTDtDb002tOkm
TBJvcw7XRWJht7CkmA3i7A4kMznNTgDP3bG3qqeQCM9LAmkSqDaeoiv23PZEnTTGYcGYWGKeuYbx
quGwwy065k+kESEVjVhAjYC0k2aKH7+fzWYNIKBtfqOnRsV3MMzAMPZyx67yvc/asDngl9uyIYQl
7K5EtxjKato4yGUkqegJPu0I8oV26oLwwKt386ydLAIxSGLd70VijHgBBaHOx6sHepNLy5ql50Qc
VMCplKe53pSPNlChigrymUC1licRrzyL2fDws2+liuOqMkpw3K3ljWo1/zTJQeVosGczMptucRMG
vUo6HOUIK294315DO13Cof5yEAJ3FTrPigs5AD9T3UOuY9dQg380UG02DiALy7N2PIJh2SCNVpVd
iKolLFqeeYnl8iBIFtLS3e7p6ZBfSNTccyURXnR5MTL8RVaPb5t1CFZ++4uvzxgYheKiDGrr9VC/
lwWeFgEZLkOFmQGbzZlI6TSLeafTsuQbaVbyXCBvOXY4n3fyBEucOdS//g4gEX7sQz5+GVQ9MiIP
KoYfpjK0fvlYL4mVKmVovmx4cfY2nYYe1VTBE5l4Q23a2t861zacNd3/BGTnW7SGOISnPfWOhJZU
Q7ztM/gwXtQ51LrscB5AUkhxHaryIc5FypPbB1QgH0aa3z1BZGR7YaJJLKgkD34I6xOKEIdL0SAS
W5lGIaGqyR/ZfRgUmI8m0NqdzRbaJpUXlB8O8nfKqLQJH85fAUJV5ybKI3TDiNH9xTbBifqb9OcN
jRsaX5VVW421Q7r5nRj11Sl20KcOYNq4oNilEoEEiw7oJtGHGqFL0Hha7uNadQh+gl/0I8yW8bV1
FwmO25y9l3s41O+ZefO24fEISvL03NgW/NBnZ53gKFVw1M0AguMLS2FZYSZ0n4qasogUI6uYDQhQ
j7Q/WeIY5Vwtgj197biHZOrorP/Ygjaj3pbHTjIJzssBhIhtIDCProuQ/O+HPNujC1Xaxzmc/C2U
cMgPxHc7VuMiOycJOZ5yK/pBs+OzwUan/XCjfdtV5LNdI/qodx5sRHK2TOW9+lmnyf2IRaxvnqTR
ki6d3nqDedIkQRt+p3kGWWbZOPWtYEXMhT4bGsAGg3woP2TfWbiCmAEbFpxCQyZVLRRZYzb3sv0G
qYK3+nw5iabDxxUU4GiVMMRHQ6g8vPJ9TM2GEK8JWBqhXG8AEly73hP2pjkKS7OAJS1S14o7xdAn
2NXvSGqco8tL+u2H9QXgKYUTEoAhJgMou0nI3IMZrm0G42UaJ/mVYZjnRz17td13XGJg5U6zykK+
/VWmuVHvjXgx8SDZ/AEeZgT0zjLaYgM1JMUvqKRirOPWLrUmjlEWg5kJs2mYGTQFUR6vKx9qeoIw
4V0p86X7Pttlj4D78kRZR+IuomJ/R+jx/IGnQUoaC9eM4gcZJl5xI7Il8Avu8wfPvg8qCdyTRx1O
VZVgkVXz5homSBYMhxo40D4fOyAzV/F0+CGlwlI/LcgEQdDYKXbvMXs604CUKTAIqwMnmlNoLkBQ
TaGet0+R9VwyWk0sYNmhtQMhfqovkr5BFgvr3kUjxubbK5dY01+FSW8B/wvtzlyT3SHNOwwikG44
79VkQ6HuiH/ffmM3ZeJ7uZJFLxDrI/QKo7Ua+IPRN6CWziXuRh20mz/S8/uRdK9PyflnoVQOMdzL
MxbPSazZQGwabvd1XTTy9HqJyGunEpGcYi0M9CZoHUfxnoHx71Kb7/qVLHc4B6OJpE447ksQrn1b
hLG75Asa3MwnabD8Duh1Qk8ycnI9nBq4U7jFiIBpEMEWNCLkqjAsd9QHe1H3FZRv8JtKHNCSBcnT
btXa19k8WETpCE7ATTs4PS+VnyffuAqNh3oy7UintJG2jhAF6zDpW4vcgxrEH/vhjieENCejZYfO
a/yM8+CT7Ik6l/GWoQYjFdSN4vFUnN384VEad8APDxSqpe7X9Jf5DkbrxpRDJD9Ho802uu50BU4Z
THUEUxONUdhl55vVpgQ83+GdvT5SW0oQK4/f6i30PPEINSoukB3fBqo+5Mxr0syZLiERO6mssIXp
ok+BaWkhGwcfP6HQ+8vTNqX5SgJU/EXiVYqNiomqsSTnJvePVqq2NhE5dNAh/1fQpnRmk2ul4kxa
cOES4Ry+FBOFzSIZtX8eu8Z4FPYnzEFWDbEXkeq7rvzVk4J/SuYR3YL3F675H2VTj/Eg3mLDOdrt
2mQnc/Abm5dB3QgrmL6n6ARkweykm8NH/CKheR0ia1DXrtpfnIr69GBhij87AwNnKpvqraYdiCU9
VY/V4DSRxveVv2lLE1eXqTpLWKSZ0A2QAEm4y7DC9JHT5bMBRfF2+54Z37WOcfvUijkEnx6MQnqC
HIgEa3Y8JNcS1xAPG+u/f/Hcu0OLgEREvhWn0YUd4Fgz+JFnDA7yjxJVkKufhQQkdMjHFkR9XzgV
JBdaQlJLt3TCcKPNmFKH6aXgMSmidx1C6ocP5DSaPQi+kGfAc49j9P3VEM+3eCl1kL5diIwVY4+O
Ek+9H2PmME6UCtzY/P4q7gg20f3uiL3ZjFJnce4IHb86cEBT/FvsxT/dY7vr8FF/V6V2kLXIkOVm
MhLfr650YClzqfrWOMMMUtzTrw4U0obXDeg0nmYYgPL8RlJXrp5Au3aREm9eE92E0lv0oV67xuOS
QurNHGj4/yvndQ5DegFhCMddhY9MTdefXmTh+L3EZ0k01khVzDHZRWWB7gwn5GF8C5jRF5QEqzU0
YByv95NIurFLFs6H3QDSCMeq4WfhnNPZg6Z4Z4QuQ7gE4k5Cw2Jd4lDLnPeK9CIZy5V6/TX5d5Te
uRZ1/VHk1+v7dj4RgxQxeSLa/fPFFCv6OVGgASZ33TsTuiuOnQICvEm2zy7oPV9mdXSMFI15osxF
Jucg9HYIjBCex2+o7vuPX5WGPaNdVmpELgNMfq5zTaFREdEmuI9rYJtn8YrZeZAeZgvrc+5k6nsj
yUD6HRg9xojuZjegq9QYgZBADgqXq9TtaXCfU8UOEpDhxn2rHCcpDd1tMnsVpabXqljthJkhbNDl
RO7v6SlHlwChWch6kIz8HuDw3l3nXE4JdMwumis1A6TOyN/Mqxp/nVfKsPnqAiOOlJzWTRpx0YqF
VZcad7jro8vgNZQy/y6asFQZsmrL7/UU4QkLayPMBxzQmOzuWu6uXal2Ljc35kh8uY/rzYMkvhR+
f9pg2eM0At1ztX4uQi2U4UWnzoJfMUjOt1XBOSu7hcvucJk38zFkA+uGygB8bTCMfDoGWW9PI1gz
gy2IkzutPo44aXoUiEy63WZHvdqxjyWBnhvmuasncpGoRuj+AlCCFHA6BSCM6ryIgqGQgv2/DuC8
QjeW+WmrpNDe6oMuuqvIlf/XeVv0Ql9y9S28lqEvIvJS+beAsneMRaOY0F+H0x0n4Ue6ApHPjLHC
99vxM3GSHLB9O5O1MWUshG8ouy47npFT/6gkJOdaXaLqAZMQfXuTbrvBXNwd3gPECvPzq25moQBk
ItejVAiAsite/MaRwyQOuOFySu+wD/yWsTtiWIJ+3JYDnzhEhfb3scHjiNQFJAkcSAGDcLc+/Q4t
B9A/2wlKZ9fJVw4MeyPF//g8k+ojBrfJOZflH6936x5iAH084IdzLwHXhPjwzPIqDma3PImafhmb
ibv6bEpta8cgIK5SJ5dHq2vHD22zkNzz5dzGWscwcEpxaLBGHh+JpP1fZz52w+y9sb4imtvzen4m
BkvK1GuwXcV9DbVFAruDs/JQJ0pUIRc8++7TQX68KB5GylSbkg6UxqSBzdal3KBIyoFaa8UqDbh/
GTdiFN3q7QS2eaj0ug6eF4Z1Du2+0gPuK39mDAWEugrJQ167CZl7w9AtVkFISCyH2gL2WJZMYzNc
mLzfyARfVuXLh33o8yE3zAjkrAA2obIOEQUd/TpgLalxx7Zl1YDS3OwWaqmttSVek6IfLIPtUSsx
C3kkg2D1Iz7DjY6FVbVli8GtQNPlvlLyuKWHNpjhRofOxumv7/Qwj4emcdUN7ki7Sfi0p4mK9g8w
/K3n4ZB4diVq6bLxMAAnSBhHnX0q2cwuvne8+2Hz3N2Lks1zKtok7jdIaM3/K3qsyyEglhOWY8s2
EZw2GHNhuyp69pdkknkijyIS7cNG/MKDM75U9uoaX19WrMHPhcYLft51h6rXUE9qvMptiFPAAsCC
Ophfb9nNNWnJwdHeGcWVYfIbUcP/2DxnifC72VsaXzRm8Sy9aziZnbMO7wpX+wk5JhxyBcEraC0Q
l5jzP/zWxYFIQeIcc6JY6Xv5ZuIwjFO6V+ClTUjETYPNjdH6qxY02he8foEjtbzc+iqI3CChBLDN
pdlUIoXxYS5iKYFeD5U5/T31Ff0nDhF9iRVbM82AOc0KgNBXBnvrJECm3NlaDN8OgS0Zlx3L8hDI
arXd4bAr36DLTdv0gzgdzuX04Ozc4kN8STd5J4wITLjZzwF6Wk1laecj67SlfycI31lFLHQN6BSN
nHAR+xOEfu98lMgBjxjcUDjZElqqmKVh9IiuUuwFMbWm2UIauanLNvPZNR+b3mhMRYqdPK7TJA9G
YLERW+GFbSjrHiJiTxhQwFzN1ZpzDa+trJDx2nSPqpenuVTou39eErjfSJFmuwCC6qEkCXe+obA+
lMidHiPAcGj7aAh0NUsqUpH8rxpQ4giRMd/bNSLP/Sz9fP12UxBejuhx1qMuWGP6v4fNUznHYuaj
hlPy6R/EsEgk2TSQ4V/YSDj5ffTVU01XB1DoT5H8nX91cxnWjr22C//eSycuHTbO53ZgMiAlIQ5V
LZUiotdoKd2FNnqbH3vvpU39ymFreahNIOs6zEOuEkYO2O64gFl1DAZcKymkiBchMSKV8Cz4+ELW
A4gMOOlMkdk3TtwiQY1dz/HJ02ClhBBlb1+v3cfUmErCUSZg6rofyejMJ7sn/8tsqTJ7gS5h4uHe
9FvjiXmGgK30zk8dva7cZ4ovzOGIaZUrfehm9Yrb4VZ0VHm2Qpdd4qIeTEmMRBq2aEDBI212sz+F
0C2a6arwcm7Unjtht8XcWXOekKUivu2N4lKRxxfDILJbdugKYDfrKgDhpikdSNWrroWeSdORNyzP
tGU564JHN2u1JxJU8iEIzP3YTttRih26gspzqN+TBSr4rJNLQ5T7eAaS1adaYM04GoU+/6WNPn2e
p/cOM6BWHSjcusb80NAxNWdYdwuOp/txNrykCFwVi/WNH0nGRQy4jziazWYhGfAUKGnK9s4afazG
gal+A+lb0jhp0dkPnajuWF+V0m6jq5xqX+/xCl33W2RELXkkMybWPw/nlHH/EE2b/VwdmAxBeNVS
bGFv3lzuO1tanu4n85SXYnDDEyv2bIkM4IeLsrtA9P0ffWNnwQTfT3xBQ87zB//yHbW4td3SAmo5
CJ0K3rBw5gL62qIHFQKx5RG+J8pyVqtQ/eTv911E9LgCv3yBSgNnI4mfVGxEjXZnzq/hmZj1rZ9w
wVsTOC+IpWDdGhwEOtA90KhpTmRwd4gDspUqw7iOBM+fxHByK2HWZicVpoXADKzcjWdtOJCZZ7pL
2pyKhexHHiTG64EgX9+fwCJlUSv0DukcdRq2PvueLov7UDLJP4CqIP3YMKGKF5foYlfEfuXHf3be
QuDcck0uJz089mIHmNM3zB7mITjO22bwa+/osj4Lq76dvE73V/3uDc7UApFn7ouPAFq9uTOsqxnh
7AGr4GhgxEf6DAfPsLBxJxvEzPfoKYjvP/NrqlVNdKnyfHW84nid3zkIdrhYdjVAShPKQc3HKNN7
e6yeuindMSAHdwkcqxR20yL8C2qbu9wP3A7jd4IlSlSOBznhBVQYPKLTJJT5hC0PV1Em1BLuqVUP
BTI22mE/qBs3znwaZqkrHXgmRdKWDyh9DmPRmuh/EsqarLv0ii5wJlIiSdx67sRAc132a0J/chIl
HdNK/RBWQQ+kVhXnNlR0RfoEr5ghY9osXcU/56PbiHB5PZi6vT3EEHWqUBWI7NfdayEsKGE2ZHw4
gH4sLOou0y7tIx1JwhXdKwXq2LW2cwphonvvbd2G3vEH2cDF8UVhhaahR3iMXfktw/FRX9ean5Ek
tFjkoxuk52lXtHjXsLitiktuTzOAHTizkc7/BegsHRcUHHtAp4XCoc4nBs3/YllsQoRBvzG+cK2M
Qr0eZRh8okWMG2BGrDjnx+9yWuoY/nBmTJX8hoKuzBI9/vUlI72bYxwZohUnsI+jCC1/JxYxzYYv
sTREpKoYCl6+H462/kH0+g4NnZV6+ra1U+rqhbzEGi/yC1J1UZykSsaIFginwCYC0LCPedM1L+Lv
0eD0OT1IdgLCN/oD51IyUBJdTMVU5HKDS1ZzwpbFWBuw+pGyN0qovXwqGox9ZN1yndut0p0RATvA
Yk0Bz/qJOV2op1RLBPhiVqUW7/sUQXknCj+aGxSPQtqJ8CbKGeVO+n64t+Ty/1VZBytpzbYEWWH+
O8uHAHSHvyq9SZNQ6xRHIfaHeMvP4cq1ty/KquiZSsMUyprX/0W+GRzAdHJT1uMhpBvnJkJ26lKR
QR7NyunIApCTZhcZqcZ35uAvA1RMQZT2+JAWy2sHMja2RbI5JfCGrJ2nrqmbxFdrgaH51+wISD9k
8aJQKD/ir/eNxXDnbbN7YzEbdOksM2EspiXgH9dLs18ZYEIzxSDohkJrA7qZJhxdNZW1N3ezdlAn
4H1RoaAN8Q0cWRZlg5nVdd2leijkdgzg5bLAhWFnt/n5LnYuEWJa1GrZLHhrmg50I3iXfcEA1w9o
fRc+9mCuqpPe71aEaYHqIblnhI45O//BUdh6Vf2m4ERLNsZF57p+ujplrDo0+pDJFSwH59A7YZv8
6xaFpkbVdCj7WlFYUTrT0PoL5JO9n/zyR9Bc6xOyvtffkgLQSRpfP+FZID/S2MLCvEtDegelUwTl
dy/RDgjNItXVsx/dmRPA6svm51you+ag+CvchNWCNc0LNZRbEzKH9Cs2QVlPOTH3x6sbqDuY3WaM
XJuW74SD/gBdGIopMyl7nPfSk/JBd2YlSDG8Jv+EN3V65Eowe4YTTHe5aVEqJ1VKkaHnDtZ4PGqv
LZ+XqhcPwOmxLHE+K9ufKkA5NuXP72mtqLwROtuqb6ehUmPjrklj49T+vMqmAUC1qG33jAol3g7r
dTuayt3KXVjuCzpzptMs+VWi3JEd4SJMn/QcxNA97yAecZRQXUyKGt2oul0uhg/33xtKRYdqov+4
b1G8QsFtkrDGpISwQJCGx9pfxmU1Z3X4vigPOAXgy8WGEFFrJfKlM3WngqG38p4pY20CnTne0Y5q
43Q+e85lPiMpw7vn1wJYK2zpPSPZNPcqqkZTDLBsga/l/c5uZM5ta7DfuGvGFifhJZ2s+DhCdLdV
fXWgxSa0fDGgyuJT9S5gquRjhxCAhnAZhDScEQKTNQQHhfQGrmcceY1pYZ7PHeGer80uFeASyBMN
tk3WS8h0kSN9bxotjCYF0CggHhYbrkZLVNB4PFD3YpTvFniGk4RLh/nKry2w1M36SVQKFhqW5alP
eRiUIjUkUQqFyfhDdPDmsTmh/I1SbegZP/Efs/7k3tiUZz3KFoQFTd+8PlHxsUkcGp80SBzQy8Pn
EswchJBPnaTpx4EfN61iqQQdU+VfdXnpfH+1S7SSA5mGlOA0Ph6q3AIljMuDG+A6Oy6pX83YVzgn
aZYL7nvNYnV4j81/6vuF8Zy3ZGKVe1OtCQq2cgiAkkB/SC/a28L4hQ0RYvwVoKHi+rAhKobPgLZT
Q1wGIORV+i1RGXk3ASaf0LOJwUjpRjb2UfnLadTxVStd+6TjYiD1zAEPVvc+h3z12dtTWwzeR9+p
FJiqKsMOKMIskm8HdBHrBqEXUFPnxkLsex5v0Z0gqnIVuiB5rUCZu6GCI5kIzjjeD2ia4BtJsgiS
RpfSed/pf24IiqLLLqyJwSs5y8N6PwzNg/foUis83WcVgL+ClHIDBAYgdnh4RhnaNLaixHFsUfp9
wI1ziTnOAznT/Uyt9xQ8GLrqRCODB7l1sPU+lhEnNOyFYqO0n36zeW8A3dMgxyCg5FTWVmXZCcC7
NCACCId0x+nSLszHFxO3ppkJn0dWlXp/EgtGdYSNTVJ7E1Mc9P6amrqMKasvr5vLo6Fw2kQPgVnv
AU7OrSbKwDuz8Sqi7AMly9o/a6/n+DQVOZ7cVMNo4KAgI+yLnY2HvhIKl4VOM75+NbIJcntCza6Z
Q83E5MHdAHPrm4w1ScktLXP2TZneOq1F16silkHQwQwuiwThXmE0LY5i8H4lBSplj9mG0Kss4+H7
1RS43JhvSkInaCqXLVRiDrajOO2WKhnVHkg2FkEZZInpFYGgt5vWPDjuVLJzbwN6xclGt0ktA3eB
QjIHChw68T0em2ED+/yo67dnFOBhG8trWlGwabVY7KTexhQT1oaMwnEivs5OsemwLROmQ2dKgj7w
hqzKDh2q3IsgaxDGlSnpnOjI+6UsmlWOB+dGeCd6OhDjwDpKbi5M8aIeP3lzCR4ioRt8jHLCoVJA
1YilaIdQi3hT/zmqZnpN6DRMITGEJckwEEa7ZXB4ZnQDTHdRUx+b0BE2tKV+5CB5yQfdBskErw/9
LU8hktlqy5c5hMOhSKZ53DoNo7SGqhsj21fux3Iy9/VQVVQMQY4PItwe942/WKmpdzQtbD7m7TZF
ZH+GCh60C463TbEixi8aafsW1xK95PhinYjHquFg+Az1LequTkgX/aF47+q9e3TYQBP/0IfRbsEL
VKee5UJnRS+LflyOBgd/wshyOsHCzA/bNq9nRL7GDaX7ZQGxrU6hR5U+x6XJR8Ms9oW4PuLMtZci
qb7EOO5PE2wQp7oGD6Gxn7GRRJxu8Cyxg02hrpMNX87idCkbgz+1cQqH4OitsrwYQ2FFdCQ2UDdl
kArvvLxqUa9+8CmGNxLoRM7ngePRBIT0DjHRmLcJhU7VvVflIClIXGvduT5SjEmzQ3bapYGz8fHP
Ki+ebK+Ox4b4psX/iQG1ve7qbAD0FqYxhNkYaeR3YzqL9m0AVz4B27Msp61sbf1+L27vnyGPGRIs
C88jttn5PnIr6tkOmgZUeRWr1XYGPRPKEvwIFfAT5bGMP/dCwazws2rGK/zOJy+AB8rsMMA0TBAw
bBfDtqrFX5/PuuisfvI694CXwSySLLPzLwbtAmLdhhcDdd/pv6cY4saGr18jOhhbWNn5i3UW9LVE
USZ609hqqCGxHOhzPAYbtJl3165b+K2aL6SE3TusaIVGpradca7OkGOwzXMaEror2PEdMCSLMt/k
GmjaBs+KyYWGY5GCHFj18k0VAzABC2uhiGgjKuZc4ixDGBumgJ/Vp+SMZgB6h1jAxTz33los0kAv
pgCpnAd3fnFNzgDKpzfCICmSR7XgU5rcftQkBSaKg0+w0Bk4pAHCCPpSia4I3QYBx7ftXBH4KmZl
pyQmrGcTICZzk40pqZbnlFLWws+4vkPT64cJaZDUTfST+at+ne7E7Irc91OEW/N8zgJvS5pOI6YZ
I3gcCpsWCp5c+1Njn4zP/5FvMzIf67BJLp+03cOLhkHnEa6eSqxEekDalGujZAl4j8wvnhNcn+Dy
Ojjxrg/V+v0MiEBQo3Szkj86/xmILEaQrCYTRPcf/DpcsT2I4QmZfnbPZDkOnNoVw1GG3kDANam3
PIc0BVWiwgM+cf1iq1UOdCszrHEl4Rag5t5w0zQW+KlIbzPeTfmML4jgI3bq1/8556Sb+Dg/mVbQ
cjqQABMgycg4DncPdQxC5fmMyKXdoTdkKGnPNT2i600OEq/9B88QvruG7/tuOeWtRTG6rgLenMm+
iYeEF3AQf5vfXcre9GYoZbHVT3EmbLsQoYbnEwqNtsAQdqHqYrJXqmzAQSYWpRcIVwNUWpB2aLVy
LG8fkpq4hwaPdEAxCO9XqhSsVdkEPyqjNu18VtS3rH6h4dwtM8CmU2aYswt8DE9z8FxVPYHxdFFH
9RcdOdzPI0BDpLgMtT9nPNc/aAYm2uuLhA5EniXW7tMJ6qIpM317V066qs1LU+JzzvXGOkmbCEhQ
ecHWjZ2waJWxhERcgMjhyBI7QlRV1ZCojIDh+N413DL2rLS6cLeQVocY5OIlY/eHg4BN2z9sHFDO
5f9+Bd4r5U2O+iqbU2nYOrQc/gz3FgXQYod54CmF+zVP8WtvgJot2VDdw9ICAOH/qF1InvQ9Z5RR
F4mAjea2tYr6i6lAT2hgTVLa7iayMLxExz7+gDh7B8TjZkjEBzGzd6433g0B9xAMYNsmkhipYqSj
u2hgMOg340sgvJdhBKKUNbJv838YHOw1H9GWmEMYdfD9sPd1Kw+KR02+Y/lsP6aBQhnq/cOIkmL3
CTstV/BWxHBZipdxc4FYMT9zfHHvb6tpGoM/WKRKeK4FAzBqWkNrYOBjR+as7DYJ2ms+/mkap5XJ
DYZDIjcmUabYYuUvLywxFAsLqaWOhuNojKY1Fj4VgcSWJToqb4e3Kts9ndcjM1bgRE/VDP3JBTRS
ECFjJma9j99Z3Or7ubNwO3S0HAT6AWIHbsR80Kw74QZ9TdP1RL404xHW1sGEHXnGynmNF92/PRaX
ZA68LsbfM+oU7yNLXPKKJVX05LSOxa5oxdz7JYVhBqadDbjZwjN5vKIkQlqiAHPZs7IYnbBomhiV
WIV4nw9ttaBYquFdaIAzrirAV9dFgfoToheOQhk+5NvYFaWGyVHKeEoILBQnUPtjWCpWuI5II9rn
v2+h+09tgKvpQSAGQpuc5aW94IqAhiMlq//zBFpBeAi7iGH025g7GQ0AGJX5G/qxfQ6bOh1uZAb9
BTqSXbBSEHfAqwTgeTmtzOvM8RIjHbG8BizpHohmhLX1JFTlnyBiXg98N3AFnfNCs2jrKqlhrhVN
NeospZHGspW+EUkElJXMA5eQB4AiICw6Py77VqdZC0mxKgY/pzagmyC2y2ExY5V75TnttVVyVMJ6
xvcxzWlOL+c0hVcXTofvDokvF9vUZcMn1z1zZPy5r63zXz7euCxwGOo9c6Lb2VgyuXN/fs123brc
g81UvrWCNcOEQZY/5NOzzw71mxX+H9+No58NHNUQbZINBGWUP4VY8FXnVgeqxSOUGJh+n6aAjGFv
BNqu23s1z3KzEaGndzZHN+SdLRwrU5O/oC+oRroZVmrjmPJuBUAvpMmNh6dW5j5WH8mStAS7YGID
QZJZx/Osq+VrCIqqmblHrb5t2ZSE5eApn5yfoHbiEvQmNi0tmzimvLCjcEeufnQ+sQDtuycW0xm2
zPMlFxN6DYRry5T70VCJ66iSQFDaJ0RWi27ZMuiOmyGIZcQHIUXYRO5hPxqGT1lGQzAYLb0tsICs
mnJbMA0CyTOSVQryrChVc/dzNT/53QCx2CnxRW6QCPp/Al9yhdiKMqmQYZA8ZVeTdsvFYA4CGLuN
ThhtmD1rFXcvtHlbmBiGGsQCe49aDE39FqX9pN/F2aooeRe55qOLidD/eKOiW0OFlNjZu3i5PJwx
TIG9aSggU9eXi2UTgQcUqI9CUyZXY0X2cRWeSGEO6LrtF7dYzgJh/X0sUvdOiEQzE5HcRW402q4E
qb0VyQKdnfqhAv+vclfP6QWIUfAyJnGU6wGxI4Qn+ugmnVe/3JmphCsSBSPsbGSj9ne1xleP4tEF
MWW61zEisIaBwHHnQL5tqjeNx/LN7KHsfUqzEQDLGlQpC3uid7DNdKB3idiFY98+3XCxKoaT9uir
9ScNZw4QpmA4BjKF+iDdYI/6vPyMuaDVB/ZyBKa+sWtxCL0nm+98KrUhpt9SeHZbOnnL475VcivJ
CJCti/mfhSfSaRMoJ3h0jSVMrmVIFUqzWI6alcE61PYFjvi+wUIUsoa8AnpLg2zd24isSu80+dmR
RZ4mVUVtG97rWz1xUNWrxVD5JmUdCKqmF3Y2Or0z7fdqu8KTLeJdjP7ZgdPjKhyuLuo4XfiIz4qW
7IGSv6WUaSyNCKwDacY4pYI5nTmdAk+yg/OUqdOJKNnBupIaV5zzYjSLjWgi9ax7Zn7MrJV98SoA
cjnpLitUJBpQH6LlT58Gd1dVJAK8Z+Jrrb3kDGNXRZ9/yfi2cDToYewJHUfp8aARCxb0dzf/LJok
CnGVYCSS9Z/iKEvw+EOAuqngwW4I5/Esf/IzmEjLPceBI2VMPn/1YNkzW4K4zNgiu1vePFj/JUD1
8Nj1XpfyfiDW0U/Os9JO4JUDYZZ/u9yDuDgnNZKdjmqbtZmzZh7kgk/npBv8PCmOaK/Yg6+0JmDY
xn69uTUZkBxcvGIFX+AJPNSKH7C7zK+RnTxU4EmIfVbT7ndw6184l9yq76yaTrTFDQZWf/4m7q/Q
0Azqtt0r1a8rY056ozh7JfW9pku5b4DaiTkB3UKJGjqqepBxA2UgxQZl8mM7nxEY15A6H/2qZSfE
L18gIUKugD4CWdnFHj/qFLNz5wb9A+hmtOQN5kcHaTS5BQgqEl0/U/z60uBz8IJ9ZJBXBjaDUYwe
z+9ls9vU2Pp+rQVC6KD9IRQZAyAlpJgbEfA8t1I+zzP8T3SbeV4j05+1B9JNn6WVKwBbprL2TES2
ECrNQCBaaTq4lJNMd4gcWHOewlqWoHKljT+FY5fjhUB7D7IcFRrMMuQ6HZf+YBjrJFkB9CwZtiSl
eaEZTOfKBXFYaX1ETp6IgyHtZXGy4tqdtBR76qPPI1z28GS7SAqt0ouOC6WUZgHsQgH0PO9KSCTE
mgm8etsg7n87yB6eHR0lRynz8gRxPhcSr6Pm7SwiPjeyyFCIrJEVZU3whqF2fQ3CZDRgog+gNKts
iR6iVybGOVzTr37Ct6Jle5LjLejk5OUBXJT84906ITs1TYyOERQJO7o1JekGMvrLsVbxMEXtP4Ak
JkkUx5NUlOYG0/IHy7grTlH14CfD9JrSKwTXLlu4IwHfs5qh+XSHVZ5MFonUqXJ2eZ08XQQvh4Mw
aR2ZdVKrs+7IMNICkDMrOWuZFJfmxksc4F8AvJZjQgJrA7R9EMgjpnmB8fDZTke/nQ3TK8fCHPvL
xLCizwVzffpIQwgE2i5x3NpTmaKhguj1UQYlUzSQUhaC/3JyNDof9cJE2Zrf65OdcWHb48RB5H3P
7tAecsHTXmViiDFdr7HRoJXfrv0SpjjZleQ3cPyes9OqJ/8ZsYRxA1gqF1/zgHM89uTboc0nqLP3
w1KBNKFS10WgWNtPOVXDR4B6ftNJyBchMYXyZmXRWaY+p34eCV6EUKJSnIGn+RnVjJsiHBZaGYtN
CIlB/7/QKmH6gHqlhe8wwSOUP7WTJ3DjvYB60UWAc3GAASrY3RPX6P6fWfeduDcVWmWETgFLgnuM
FKe/oyyDlK6V494YcnPtRQlsBEISeOZkGpUC+o+6j8oDIThPTDt3YZkmKELEu+EEJAzH4gTb297U
QDxnj9+rRMtPZARzJIFgByGzvUEIHG/77FXvgCewg24p2gLFDsrShPBL8M8AKR4qQhLFzXG8mRty
E+XPIIXYeY3yip3wmhqBg1x0d1Uo/3xn5ZJw0RpxuHYlxhzzULgzzs3RaFd5IAmTgDzNEymK3loZ
ufxHeGDY+r5/nSlCrsRmyGtgdYfBVoYldsr6B2M8N1Bndqkxo3JUxze42yaP6rFWhCfOM5BveN35
OsHbD294VBmtodk0XsDV/cEmycaXmSsR8VgwazSUAw+TDU2sbqu4wR1O6jQ70GRtb5ShUH4ZZU0b
d/ha7JdMoshyhZsREO4kTZxqnhPyQLqazY1rqHct1mL6e/4VjnlAa7VxWKP9pyIudmt0sfhsDEoj
30XsqcwBAI2dviNT9eLVr8D5PTveVA2T2ILbLFWrb+TM0MFufwnQ4Ge0P73p738ZkFdzD96sj3aF
BM0+DQp829bSbnJJW8QydAYHoofD+be1aO6DqbPIMj4KwT9OmSapYHo4F3CzeI9OQKQTa3KrvHF5
+WJ0sU2CQdkCh13vL3E+kyLFpZtmijkUg5b80FR5xGVAXA/hcondHhZe2ZljMe82aAg5Ef5b89i0
iwpzQ/1FELH8Ir+CN8tB2xqJp3qPv9iutfHmsoA86Odt1Kst7TzRnU2MqdrDBCftD9EErTpldbp3
dhh5GyhPO+U582hqzvKDxhY6AR8cRF/dwKKo0TxIMOfx2nbQjJHXB47tFPk7EjIf7B/zCUMrIOp1
hUtz9iQmc75e3P/sk5pu5TWC+EA8acyhhn65Nq5xC+0LTyy3LFQ/sNPRxyEFZlJLYD/Gqy+fFY1o
e8nrvTc6mDEf7jljMCevE1iO3PyliPX3tkZBa/8Sn8fM+hVkpVMO2Ewd34cy7JMWd72lGPWMLQ9b
vRT2Bim9e8M6zGJ8uh7Gvfmjo6mBaWfwlQtxi80U9r1O9TaN4gnJ0IM6EAdMuSnFzO/u5I2b32Ji
3kEi6GIKsrfV1wwTRXsxD1hSZ4BzcqHe1DZGRwb6fQVdVHg3WUpG+HzGfnhZeixlDUWaUUg83KO4
a/QJFKJ4B4U148pgr5UyPmE/s8WUn7gsAmI0qRJ1pcYmBllmhUnEhAzdxqLQLMDUw3vgXOWzlSTs
b0lKgJzG9Oy1LJog7ri73T5KvPeUeOa/iN3ujb0Qw7fE+8eAB1Nh7QSc4ytoilhk09VBF0YC4c2y
In2xuCmqyhz1Z2WMFDi9QWVgcDqrhurkFJYeyHt0Yw6UNIU3XNELfl4XDuGmKnk+D209+Z8UatDc
NZ9SeFhsREDv08JRuYFmSsdZn3PpUkKhBRqBDTWW1rLInPQ5Fgc+DAwXd+gsf8qkGARwzYK1Sx3N
FVp6pWY29j35oSxKy3dyjrOscpPZh+Nl6QFGpa3Qq0oh4/H0IKiUfh+qY2UAqlvWwZDNRwdKOiXl
QNCQjm2ot8chB9jrjjjXfURszftdxhgamU6BNeNfye3x3+y5x6HnN2bKcF+gME29tsuh7aoLUDcY
qdmk1m7wDXaRbaYQMfltJNxnWN34yRPoB96wsyWZfKCdGdC8OnRSXpibxH8YcqN/m5597Z797Vb/
d124Ui7YBX78Wm3+x3j5eG8+nPqktRdTykP1CErfmc67r9POWsVLIKrvurJjzose95XmRAWk/zMI
con22+vNaxlE2dtJSMsjRgKkorpBX8s3B+yH/LhgUS3VXz2A3wAaOlCtqdGliQC1ZtxOkYHt5cPo
6PNXzsFL/I4oNEniLKd9SEwxgENsKi2V1tztAV4PCcH3JjG4wOVQHQhY95UmDzmv7eQJ+8nd5OEa
lGS3on6Ld9g/z+Ry4PvM8mYkS3c3lxcrCK7ttz+AdYf2LEH8sRMYIg/5txdfamTfeFBVORKQ9UXV
Pj0llu5ZGqxDB+PNIvfd7GUuTr8AVuk4OfcnE+KvST9aRF/VjVmU0AgAz6B+YItjX7JScdHH2Lz9
lmY8z56PZKdtdkcad4tRkwba9dkyr9wbm3mOKKyvZnDLSe6x8tgvwRAk5brNdphKmzH09Ga9UJRo
ZixVghxpXpjlnUCezkO1k7ftcd8KbhUX9GqhZWwcEEwtP1habCHMaLzBBzYpFpR7nJRktvOS0pFB
fNv3Us9j3JG0hRYGwVRiFAVFbyE8cQpgNap7i0nP+bnU5l3d+9dCnrymBOCPzkGgZCi2Z+BX7t13
Ok71FajvvxGSSCtAjEiPvUShoL5bitHbc9LftkORuORurgjVI15KqYlTEjecoxBjGXD7+ZBpZSp7
7UKHvl1k9gqKTGYISPWYc5wUph9+Db33AhdYlcMbjL5/EEr2SzMNS7FEuLq/wkKXKp/h6BBJBfcg
0x9/D1NSBAFQGyOBxCnwqs/Ol3Iv/UZxrPS2B2JYq/9IjkTtCaqagwCkKULduaBLh2YAWbQskZoc
8vBDZVI06qbb7PytnvCs3eofgeQ/wxxQ3nRA9X5KX4xMzANMTH4nm0PnC+4VYWpqk2GN2Pcl1qEZ
yfwX51mUlwtC7sR696plkErxWXF03mghakacl6xQLMSKMSn9rgN2zIA5+DQ0rzdOyCwczmB1MhRS
SEyX1aLlYaoR8uA8rd20TRyTEMWzG57+GhouYO6s2XpyUiFiLfIEK2oPZ3Ryru1yw7xnsOm4ideD
eba7+csditp0TYL8iW2jdHgpZvlsZq56Uann+ruqDJrTAxdJZJZFhTds4No/MXyArplpZcM1P0yX
xBLqV+U5jn3sgD9Vs6I21pgccWOTlMA5GVbnvmx2Gcd5hMWsrYx0FOah7BbhlfGmk/Od8uILMFGC
gFjavLGbdTKLkAPq2BGn8tXgPDgTBx524fqeGGK+y+NFOTzmC6qpSM0lbzbYmh8mUd+FFbOsUuW3
Y16tH4u5Ljd18vaop5kkXIgKK/ccxpTC19NKmZQVvrcfYU3cfQ4EoEcqKvXWVOaAz4newz174oQq
qi6krih+0XgNPjVYzGcfBxXvv5XTuYNFuEJXUN+CYxewOcQpyKxRNlIPiom6alLoMcxFnc8QyFE9
0wcjiqrZvD1QGQci51IL4O5U+B/W/rYjwIEVPcT+eSzC3WP25CnkQbe4mw+YOefNsBnLpc5117dp
R/UmPawYTzfUxAlqSeN/ugLEBQkGywb3ZVHO+eJlQPru3CNCQN5JHhV7eTEilLhgdXoXgCTj+U97
3kS8YFwCVeeriv2l+qFhLjaCnexaAhsUxfiqYUtxbyaoAtcLcxUdU51NSW0U/x4RSbkp5XU0BUNm
bOiTreC1o6BjtUxGlEQict72dSyHjuQ8jBekNAk4fO3grU/Xc7wV8ouVsOLiD00mFSL9j904STK8
VQB/jsJpZguPuqM9apT/QGnXbbPNAqq0T8RtWVcqd2C9G4ITs2rYXMqlLTss2GT8ppxQkvdOV2E+
4vBeVT5S8rABehjUeb62Ou48YWTeEi8ZH1b7za84AuCMaJw/TAFZ6w71o6tJoJE6UUmcBfx0fW7T
LUXA5i5qEtoUHW6KO+MWSiP3MA5u0Q8LTvdDcix5xkK2PCqyBf73zDJuL9a4b3/pWCFdL3zjjuY+
D7l+ggQCG7X+8rbVWNYRZYI2gzDFaDh9bxmaGHQWk3w/PxrCQHnm/WzmNfKtP+230Ck/dhLQ6tKT
itMeOlY+Zw8GFNoVIeIpDaUunhyK7eTVrQ6jm9tMMEGB6AM38xaJRtxOq9STbgJas3Rqg6T0FNc6
GnTTiUoPtfWkFOYHL8JafxckzDGw5cy0RTG6nkn8sfOwLOXMx5F1uIu/EzV4/zq278q/8L2YF2Pl
dMjadjtf9Qb3WIkfFqX5/8nn+xUi2nt2VGREA1Zf/im1a/LpLaNybDK8RmyxuE5chr3O6Ny3XjAH
E1jD3k/OaaLX6E0rRaXV4uLl3FD9G7iqB1kB8d5R+6wr/YXhFLInNupfPFMafGU/vXQpH+gHAZEC
ohVm581YD4NI+VqzP26T996SF6GcItUVY6GozqnaWSN9MgNpDuJOwcNAIU3wgP1Kpv783Fr+lTon
Fa/9XtweD5f09vXDj3LOFHChqOvBmbonOzQP75SL6QArfhFs20nPSsbN5vlzi45hGC0E4/I7ouyF
YnogmpdGy5hBMywD74LmIawXughhSbzSv9O8MPMps7KP8/+VBzqAo76qeNiS65Pif9e2M2cfGTCM
mM/VC5wrhqxFRgfH6SVAAH2UQ7o8DDZy0m32S8EiUmr7KkzZTDfQpTylh/VLPZB8XUK2F0pM3XXU
HfK6EDLReRPXgc3VQIFGq7XhzHL10Ww+RWTHkTSkz3h+EclYCTfFBgxTwIdYtl20Mw7PmFM/bax/
142L3ykRVcDhBORq+14gzazYy8oJN372ZEFMgjfyy63HMWm1LBqAUkFujhn3LbQCk1ttoLtusHr5
Stnj5UYwQpCVU4lMh26M2VpGi3rl4go2Z553gpp+CyZN5kuwujPmlEbkwbSjhgNlVJM+9ebcggyo
tzPgx4UMtD0uMBb/TS4E/zjpCA2h1bUUlfGbQ+juwhsS07UlHBHKVw3KajQHffNcYESBS7wrDHar
RqETLN7dx6Mm8WSloXslzvyemiBqTxyZ8O3FXEeHGoJHCtBNSk4aN72aosjA937hWIBHfTMPhXzK
fRwWoKjnj7/E6QguZK0z7ghJ8LiPTFBXsrMhgYdk4XnXZIvDyLbvyAzKJBXnnHG3kWLT1kE7iVFF
pujRx3UCGF/EACE/uyst3z3naDLkITYL+TKhferF4MMzVjLiMT4tDo/4CGFLPwFMhsnPTGya7JbC
yYVD/+GGgehGFMBq5FvSWp2/3Z+u0pQBQ7BVnTAyC2dvCIccN0vKXJciJNLoX8/c0Lkercumzvoh
uFfZN8CPXqXe3M8GL8X/5ittSLK0aXIB3JLcI3kwLIZ6FJ0TTE+JoOuVwJ6rG5mp/gWXWXZ6UnkA
zwpHTyQPM+eeSkiiqaKFyJOTqZncEfmSzjTW36ORRtpNXkEsZR3jjXFZ3Cq43kUgjtsK2nUsDU2V
6igWxPxwKQnlTyhK8+nn8XfdXWS9J4d2Sf1E8O6M7RklTXNAtVH7xfMMX6y+mTlfen5wfqZ0qzhi
5aeRFcj6Kt894U+KYrueoeQL2D8zi4dPi5FbsU325xxr3Y8sqOLJuubfQfVbunj80KLJ+Ng1jihl
VY35Nhg/Gn6awgPlmi26Q5DXN9HyxdFA1S32YdVdkg7JA/53mZ8MDJq4Swia2cbtXiy/xF34vwBv
VBgOoCspyZGx5yHnZFxbq7ss64RrfXWJvDydshbaEpE4qcKZccdaz2i0tWB0yz496Cy1ymhZRLgK
WqvOPjMRemgSYbR5ii2GEYydENf1bVGShjkSIviREawRGmsTqGiiLGvcDWOLGtb2Chn5URPlf1F4
jQTUU3C4N4CoRzZpW1LKogaliARUfhuaLD7MvSUJaolNsa0vbSUzgF2yLpCf5bn6SxCELxRzxpDE
2Tu8zYEaI0a6dEy3ztTciwRQBWuBoLeqtQYyAhlVviuZKRIULZRhrDfMPqcNkNf3Q/m/4o3yvqq2
Of5bySVv8EmwGhd8zkx+QbF0MaNUqa8W6xlKnzWqO1UUNE8sruDAkOzoSjSVfSD9ci887Qq77tnt
NpPDZh5YOaV/MvqTIgOGLzd0qe1P9VsACWhiiGvF6XuX9oSzzTKkbzQpS9MhhJol0u37UbiHkQgs
KNI7h+2lz50eePWC8xfl4Zua/rrwG+CL6GlbJ13lrhxQwvLSz8KXLJwttY/h6mSAfK0izHJaAkrS
MSUPP540gsYBHsHcTLSsVxV6syR+DcNd3t9602SC9FnBFyfUxShvqKEf9t2PAjKVLCa7qe6etEOd
DvHze+wyPT4BznESYUhVp7jcf53WS+rWu+ZBM8SFYuikYMnqaFlwU9j11G5v7zYh7f/Zp7TcxaIY
RxyHM5zuVFOLrSYsQInr2vclgwOsNTk2IvNb4k/YZqzELjAYOvQCwNht+MvP/gUM6Hpq0Fv2EqKT
5s5ANsNd1Xl4A/iGP0S5Oz4NVjPBwAF/F17s00d51bV8AKwOBqR3eAkvsyB46uxx8eegjnWf7vhy
FRjChShyU5rL8g5bekEj1fpNgghNDbQrVeTwX9tWkxk94h7rH0dlJUZZGKPWLl2tCd6P7yhg2qzl
pxhMmDo2h3HmUkiJlvjUbxvSaaeElOSY+WQ/RyBQxo8XzSOTv93RkkkFQRUQuEo4++51eSAXgDqe
ZVETFhGltPmmcKS8dg7ZuP3D+SEGhI+BfmMrWnN1iHFynHv8eyWXOn8F3f2UDvupADt+AFslJbo3
t3xhJBCWQ/5zG/qvYKkt0xl9uzQcEKbM4BbPg+mMiM4N9j21FQkXttpTgm4Lzz6sE+AAd/Wu3cqe
iTgP+u1UeLqJ744tMh9u0sS7LUBkwiodJ5BY9Y+M97c6oDxWNNtD1DAOqZqfWaXhAdpDGiq1oJDn
qxEmD0HB+TkyExNV1dvqd6fFqcqWe3vNq7IwFv0J487vlyRoNtEjQhNYDbQEIM2N/lCMAd9bcJbM
1apb4NUQBmA6uhEe4c13ihGePh3PGuh2WA88dROfk3vZa0PUfk9xtxiacb3vZkiT5SyHKCD0hrrl
fZKjYbxuDB/3q0fX3a4yrK7DATrOyJJh33wlDRdz77PgUWYwDSZ87jfWuu+syiuAu1KRslWiJd74
ynqSVxatJNKDjdyjFifUB3ixg1CioQUhjy5d77weEkf9y9Fb583+gmVbehuXvz27jr9VkR5HqNU0
Gs5Y+zRuBhwvBjQYjvY4SglAqvKZsUyrToOGMz+NG+jrGdjDjussjT3hlhT9pedmMdV/E+3C+qxR
2zHVSjGhaXYjaCkTzu7z3KTN+YDUjynOHSpfuu/1cHgftCFcRtm71ZWSMPAXJYMxi712qKL/Jhri
DbPyjfcAy+GLiEGMjLh+XopS/97pkADwgwj/+TzxKhCTmqiqmAizK5QQE82Dnvc5NoH+MNSy0UnX
PXQdPjf+H6OugGpF8BPrapQUCQhib8A5jQwc3GPfGWvAg1VfggfnIzLh3RTs1BBM7YMzkmcJCmPW
5qpghklSDrLBAwfOjOlLGHwnanystEMoe+6N65/CNl67g1u7Ro6iczZejAct61/TWhESeDrZScke
41nPUur9ej/U7EQhJ0OADUmj4L9S9du52PPfsQIoXqw90LFWJ0hPa4OLcUyb3mKyar6h+9ZHbfuj
tknn3cMtcTeosCzJBtsbvxXSm6TTCMF3GlgN91Hn6i4+a9apt+cAHUXitVhq89yLu8T6sATIcExp
qdvXoBBrcQr2PagZjjzM0RdgBQRAKqZbnUrFpcG9WJuytOp7K8y8XFPlLDx56w66ICPy5XS2Jd0T
xgsgx0SjkCwxBcltj7rA8MBGUYA9xwAWK1rEK8tp/4OwIw0Y4XM0xvGTBK4/GteqUukTu+pOcVvi
ZMP5/Y9yO/gvVu/MUKe3TK6Y8ngvnjSwN1Rlm499LS/kpdJ/2ppJzyDlWQruyEvEZZX/GUqRwiw8
d+eDEglqIi6oGjHspq1xyfyFNuur6+9Z4LSh1QuBhk2EREUtVdLUZ0G88rB9wXyEX1V4s8/K6w39
z2nDCLiGBCVXFkqE7sXt39JsVuN029gzZ6AEypz6s6cyOIbbuhDY2nH1zXzgWjSyfE/yFXzlDXOt
yRlCARq5syhLMZ06JSOSBIbWNJkL3MpMkeCt+flpRXfZnL+ohv5icqwsY6q7DSEwA+cC/YcnWVJ2
01KFAfp6W4Ga9teE6M6d2c+J8doRoX8v1h7YEvYV5C0m1z9PGWZHlTfYjDnKZmm+Re3lxBOO1DHE
ENz829n3G1zFlmdXoIpq8HFUYf6JSxVzoTe+Cw0rBZXPlGSZ5Mfr/z90ljUlAsAeZc3COpXHgDAc
bi6ANeG/25u7JQ0hQPSVioMClClj24jb9hpuXqTeceW7v1HpHhUshx5tD3XxQ5tWTsiif+wHlqff
QhVrj4rtyHeXkLsBycURP2blwql/iOajxuq6pnDjxv/AzGDrBwZa1hfFeaehZWNXh56zswI9w0Sn
x+qPqlgwpPMqQRSTcMH14sEOqW3Cj9gx4rCzzJhBLBKlj2HCxFzEtCZKyCy4SOk3qiahruSXt/vj
2C4hdvy71fd5cYlYPg2hoFZ2QOXdrfC+Ce3Ib7B0G1lVFKXYIQg4kTNZ0bjG7mE5dcmjnrj2VCJL
uG8CEvR3nBxmAKX5GP0EMVSHfYn3E7kxTxqRPeKrPafwRdeQ5bmQuWXZXvvucKahiDDf6JiFxe++
2TkIP2Lm+UBoeCmH5aX38YCnBLojS9KBhkaAETP98Bf6E3zUUNs4784hARgTj40hvg78NrkIswbC
No4bMlA6YjaHWafCYDwQTnIQJcCsRjhOAN0r7in/mwE+bpFwBYCzPFwuqkQEqNJpeZ6Bihk2HE0k
w8yCHmUdnhOYadwfCefBmDurvvTF7FFNcjIzoy2RQk1cubNo7AdiRrwgrou+N5NIMgnfop2KzI3d
qbM61suvF7NO/KasW8ldYi1Gwa5BHBkXCnKZVxoov+QrbeYdK+apadiF+7vi6or4+bprdX0/Lp94
jqy6ggt+u2CQeHGiFvOT6foo9kbR4ddDkRSvNLc8wHyURQP5BGUwUvZPeq3q+VPPvaByfwdg6tAR
v2FLCpw0Y7xGPxkVBtiP908/Pq7reLJEf5DZKf73KIgFqoD6WCCwjxQVMtJmqJRM6LiyTb6DJkvN
hGSrZDSK1Wi/k8tzVyuy2aIS6DgKHie5shqICOGEvMrxRVJWNwAwkE2LbzVEqCJf72eLgONl8qGh
UCi3z0zkvANozTCriTlxNq75ipK0NOGLg3paL94zRM9KHf09gmTHX4Tx2rGk3YZnXVU5lDyJym5I
oWSYIelGHNKhEJmdJ3GKthrJuy6vmF9Z2J9xeyy8A9UZA81YOjzr7b9VputbCIh7L4EMhex762XN
5mDdwJY91nejXt0ytubDK7Wref4e+02ZZ1AiYdCS9oGxmXkIwrQt6OWUJN7FSZOfMlWd87kCb3x9
cigS8ZqR57oC4rncDxjEbYYO3oVQiFXz4haPfK9xdgXJvNLQ18jdWqY+F6oxNsh+oQMLbwuoTvHq
Z/Nl2T2edMkMSHXP1Cs5W20DT9qP25VtLqkQUQlcwqFnNYarthCpcDaGcKhr3Iid5jIxrtTPQyjB
3ao8XrUTq7RW0W6vSFfKfCLZ6efS2R8o6uX31PhBEM7iKBGGQ0H59a3b6ASK1E1gy3MWyeARAYIT
m3vKvqH7J1c2BkvkoHWnPHDQzp/xhAg72u9aCRlvTGGTs7u4oOVriocIMnJ2z96jXNNgkcNgWvDu
Gm8+x+4A2tpV8mBQczqW7zFY1EbUJetSN1RTmsVp41anl5IvXP9zCZb7WqeWChSNpvtcb06p3gZy
KVDV2tWCLllzxmzPJ6eYjzFc71UqcFWXqDjtvdxa5wfeXZ1fWqrJe2z7BRb6wyFT3RmWDCFL/Brw
EmoxYMv+wddIvvwcLRdcHCOk6V6IKlm+WB6301TSi8jIMQWiundWRjrvgIWPhNM48NTxWGKrRmqj
vP5TzAJma4lmNmelQkOYxLvh+QU/T3xQ3DckibxgcpqETFrIdKP4Ld/y+COKolXN+kpBm7Z7658D
Fl5Gdk1fzW1rJW8AiTxTza6/2srpPj9WSERmzIIBgtuaMSnrdGuA1DZZxN4fev1n/iMsl4FU7wt0
pv7zUs4rp91b3GBr8CAyW5ME7UM1g+H54CUUNceMLLA3d2cI5Sy/ILzvbE+DSdKnw92St0tzxZ/t
aBoBRyrgXVR6CxVCQ7RfzCNmvc+NtMPDLuJawjRqkAu2Gug2mqHBark1kd9pvdyTMCBuydfdidRj
dTFlwpMALwa3IrjruMfd7MdKMeOGo/YXntl4SMalOTKGJ9BjMxw0Alt9uIUOcG6Bml78RneiOnc/
I36nvJRypu/8EFdcrtxEb9b8PIxEW1SvK6S/68YV7b12we5XdX7HAswbGxhWfatUZmr8ONPQ6wmP
lqP5Z028mqntOQSK8//tiHusYIxmuS0LkARKY6w56vi+8cF2BVgPKtOANTpbscwShs66qbR0rgG/
QL7w7iveu5XzdFgQ1OyJdp2th3xMKGjTrHuUuoOAYooyszSEaRj9o3PcGthZYXKH3I6VcIxCfAlJ
RaZ1DqFKCE/UMArXflgkM4r51aqZn9zClrjQS3r80XY2ZOub2HbK2qhMKgXGet5yIEcu5eVTlSTN
I0FNidEc6PcOqQRfK9v0aX4T3m9xRmjK8uWiZp2LIGkYmm1zddHH0IDSzlAS89tY61A9wd261x1Z
JNezIWCpMc4RtEJtbHAnvLZoHt8GX41gfc0RC8QcM/If73fkCf3GVcGm9JLvDmdrKA9+GMPzPLgM
RDaDueGkk6d4ZLd85uc8Yqa9I79bV1bww31Fejzb6fRZv62UeGoHNFB4atSxFxG38a141Gtt5Xll
y2bm0T9qXYpbhHOLjvNOh94H67YMqYp+7EfOpbpHvEmDWDErpx/99zYD8xvPpytXzv2w1tflkUiT
Utsl+/YscZzRk7kTX7ZOVOCBAPJ3MWHvcyBZJ7TZteFcy6vS/YOx5y+xQdN+XTPMopBpXT7EvSkP
+6ZX3Grw9K/Y6E5lFSuhs/gqL8kAOeapKglst1SLftXZcu9S/+oQQIxmqvVEER5HOrMAm+LCgpXF
RMXt5Jo+5yT4b7pTp5+HmcmXtyKj8FEB9I1hT3sGii2Uvvnhl9L2XM2HwpCe3W5yEpnQWWIOl+w6
vkYOqMYY3CqOUW5mKXHQHsw4JR7xVSoeyV+HV9xWa46NtX3I/EsdizL+ZErrE1evgAxRvb4QBLGI
E5R0npOzZzTZ45gZ4CQ+TX4xUDVNJSg2UiNvy5OWY5Ls3TjWVjd80PFsLYRPpIU5lW7IDmF5OqUU
YC/Sb0quVkFD+oMPh6m+TmKgZpXfDdlt4Vd6Y9j9J4KZ7os9saamFqUg2IkJX0B9YAM3FTr32lCs
sZkst3oEQwEsCRvdk3o89XfRxHkH2uVH0FSovi5odGnQ26wYtxL3kx4wa0ns1WJJfSs5k24lv5Jc
ofggAveO6avp6JX69HD07Y4RR70/CDyAW/XbZvLZL6+Td4S1rqP5DqWU8FiG0bn0Ae1pTs1PXfKF
galcb00ZbZkpwCNV2u7f56KEG4xmMuhJcxHjnDWrG4zNnL+7FnwTbcjgGPCpISTk0eHd2eVIBHaE
VLRl+8jBaifa41le7MPM0BH1wkf85lPu6jNsYGrIQJiN6YEMJBHiszzT4B9YqRnqGIrpsstjh/+X
Cd5713Mi7i44k+SxX4uLb/38EV+YxI1eRYHrM1fPKeZfTuf47KeT953nfVPPrJvuwy+yuLEox4iC
HF0FHlPRHxnzR9BsWnxVgTj/Y9XbuGOzUDbW0wBEjqwGcnig1zPc07BZOFGJKG0QnsAa2KcHNjpR
mKS1rQEqI62GWCkORcL/LCrMY/nqXZl8aYmRN2z1M2k0hLJRxIjoBFBKL3zHQegqrkWoPJs+pu1O
3IxCkiee/HHQwaThITsYMCFxLWfFz2zfSl3MfiywYvA+r1D9LLfIE0GGQ3GKAx4ibuATWtZzxysH
2G34B9LxXtYQQoJIxULgnDMsDJiIVPb/P7m8BiY3wVJMfKLX0P9VxBfNQDwPlS9KT5llMdDyiEgi
B1WO9GqZrW1GewLkUsPXCOA/jvx6zojY7xBRj9maq34MHyUYvA+XpjNNFqRP9eXFLbNG7IHMxgxx
oxZ3SRJK3WezMoYBh3YH+IeMUgbzDf5EwZNxA2ySkVJbMaTVZhL3JJIeW4M2xM7K72P+UcPA86kA
6AIUbIl9MaDxkyzc4BitW/OY83TojaO4xwZQo2QW2Z1FpWOt/nspjA1KUPXhlH3ahXM+fClAE0Ls
4Wp+UbWrj0T9tRlfTJUviDxw+TDmJRbxNi3JQp3Dj8hN1pjJaY0QuuZwsvhObx+uKeamvy+7D3PL
lgFm602yckA+YQV/oRIQfVaeBPLStQV4OcT0LSaE/q5ZKBEW7agqOwUOFPlTWnxOvu0vtGU+rx1a
PSG51xq+uZkH/7/UyOHsfMJjbH5mLHlhStUWh5MTJRXWC8ipZ7A3o1wB1QtBZVZ6J+gHxbVZuVuN
/hmyaBN9jiks4ifH2xxRovQp0wgee79985tgbw++X/R92QvSlccAjVFmfI2ZeC0Sg7DYYTGf6xRm
+xLjMQdah/h1NVZwVZLx3ZQHcDx2vRqFs6RzvLVr2kf+npcWjPoS0fZOFTkS9tNI05vxe8gOKGcI
s5+TY/6FP6aRjgPfhKeiieVWM9vc6BFVp2ftemOJyCPCWfrDA/UmJKt5YgLWmJKe6lR7PeBvp28V
wavl9xvkgAaSZkmGzC+FnUvgNhEbzTBDc1j/KKNop+SFFTWZq04lpdxl2CSoZatffUgcDch1Mt1S
1PZubG9tL5g8fl8iH0gftl1gOsmmSVKSEmaFNbaRS7keNIq8AZk0iIx6rlP2GrmDf5dFvBf15ERu
Vks0iQHzufQt7BI1FrczOW9yPB+BmLcmx5V/zLSzkZZlPHp/Tqfh5od3N1T6gsE5EuqCKPJL/T8F
LfKK4Ox1T/FddB1UZf3FyvZeex+uPYM+c0v9AWq5tH21RIv7vhqlmFpUnZrrKkEAb6X4vjjfZ5H7
18YdTdHeixWyiKAo6gNRP0/uro7Yk/EzUY24oCThWU7cht9YzkLrazmYCKLbDtUTWH2+fFl1Cqzk
1G9iBNbpKgqabY9HDog3w+GE5bAwu2aIRxwnM6LcrkrqHuFMN1TsVcAtNpb7wH8Iy47xWAUJvddB
3iN+rE9KKgw/TlbDsdhLhL06TqiChUnYwhLC6OlTiv9Oyz8fWRhRufow5B3DfIZfx4CkK2eXAooy
CdH+ch2khuGqvp2iDW30KQwkifWQQxVNX/2Nxs32twiiqbGwIy4eHhwwqebA0HscdJuEN4EuqWAE
BHONTLb9l/roCDYsvRwe6vbUPAFjoL9jqI+5CJz56TP990Tk7vQPa2iFfLqsWh5w4v3+eViwvQmI
lhX0Z5YQWj6W2B4royIASV3FMOqbqKk7n3l09y2TgGKfQfI6Yon855LFH+NWwBLPyxtTx/YjAphg
3okGl6yQSKVZyVKPLydxsQvakB3v+ddmRJlzxiRgJvzcRxScmDKc/+3R+PDC3b+weBzzz8R7fokt
sOCTrSDzp4suMJCSFp2UK8Kb1V85oyuOmpjK9rRuFySc82DOobP0PAPPV1KkB4nI37YijFZrWVoI
Jouwz5KD93NtjXfZP4HQqY2l3bpY/ST57d6bCiWGnU9pU7S3gay6XQMTFua/Z+DuwNMwI4AErzKt
DGydUKvrLsxjFeegyhLtNrhHuqfv5BmnoLby27vOtiArPJgiInVigrTgC1XDD0GMdF5biYFhivdn
EXv1uQJlnEpFKiznwh4E55LhVZ67K5bUUOZhAw63wQzdYIJeKu2tH6OxboDL44hQ2nGEHUkcGuc2
ki/WBxdt6On+cbEWSE2c2c0CfC0lV59A9SUX2PMYrpyIQQqQPqYWx0lvXS0WIck4NyIOllHgFbRH
o9FIP6s14kJzedz9FdCTSFpBTJV4AjnELJXEUFbeCZDJDE+N7n0rPCXlTHZ/b5EYoYFiOuOgtaBq
D+OPgWaMnwGxAD2yM+PISjt6NSC6kz9+RrmgaLaE9hH81cRQPNU30xmjHuuAsRNBs2IqqQ0hyqBa
pDK73WFB1jmpRmbJoiIMQju29BUZAzZwns4z04xB9sAtxnqvnQHH/ZQ6v3XmuR86sCDrSrJKagrz
zP5wpU7xQAgiw2Pw5/x2Q+RXRi4mmCntt/vreederKKk9AHGHFs5rx0YmbHJzZqT7egiDaI+RKa3
s1J6gv0O+H36VZFTKVlN4L39JmhixYOGql30+ssClwiOXLyBeSy+8KehcyzzBNDLCW53yKYIym8Q
WQqCk2sDl3WXowHbRflv3Wp8m6KXyGEsno5FLTVIiXs/s+dq7zKUq6izzFPsWAl4fenvwWsNyzDd
9SNSBn58Q70CXByLzKCdQon8mAbq2/+tUlKO7HdGSo563BZC0kqsiBUDQOeqQ5Z3br8TdwyaTNiB
x7AU/Z7FZ7TIWEwPbvdEQVWWbtQUyvaDsT6Ogz26FCf5qZ+dNXVxVaOaHmbmEqactq2WLqlG/E5s
NTIqsrh/w/zHCDwCBVvgOLDPSR7fxiGY/8UOaegQOH+XMTRcs3nnoA7Ww5FXSKAKNl7ZsLqQ9JC0
YTum7qfEB0b3XZg5UeADJOtnm9B+yMV5ojRtGR69TiPreeSFLH3ZlGq36euZ0UikBzFNkv9zFhRj
rBpwCJCEpmHSIZga9xowTAZ/qWbwHIMRE1bB6AS5fzsPtxqALQ8vpwtdnrOSxPNYSR1nawi9m7k8
fr13ugtg10ku4H+7tUURtRESTO50Q0h2f3S2YYh5L7FfNLapsT1pGXCtwjbRtiYAQ/5+dC/tBqbC
nCpyFKvV0pbd6rjgRBkOECi4y3w1pjmznpllf2/0+ksFI7enpqNVNZtd7G7SMeRVzxNqNDYflRzJ
GhhTdxHWCcOH+eqtxWrBBoFChEUyPgoovk4YxpgeJNkNPsilUc4BAaqKDWpo5dvKHdXYOUcvDEOM
dljiC14vBLpGzzwAFwWtBb+Q93vn2xEP4iBB85Y3wOctT/iLlNOmr3iTxv/JK+1Md1B1Za/bMMIj
bj8bbBQZfdFIi2pQ0EOJT3l9CiQKtL6Xp6a/5K0zL39ux8aBKzQzSuCQV4mwH2SG3bjuhulm5M//
Xlqur0RGO86BGkIwBDgEzCB6/lNPH8GLPkmKUwV+Gc6qnDrkbV7TUdTGnOHBTTMcmHhCYITZW6S+
BpGrKpeGxuFNNGrF0AgwHeWDRwscCX+O9a7dzKNWZpxcGfA9gsUdzeJUW89AFvpH8bwt3aQFqBrj
Z6D3aptKs1aeBWFA/jflQgfOx/EK4OY5P+FtalAbpf7aJSRzjYjwJfTWZPTovj+fMwz56FbrIORr
Jcs3nt8mx1wMMReOXEKPgVcuuAGgugbGWowWQMMEy7diLWyjxXGd0IeKyhwKeTSfglQePF7vp44c
SL0khSk2W3cRVd9WUx8n6Wm+/3omD2CKukXYkkuI8ujb1kCk+a5tsE1/0KgJ9CVLeJielGH9b+h7
Q4lDwQeAG0pV2RgCOO+SO8F21CbTX5rgbuvr3et5jWhj0qNV9/UTAgQiZiKk4/oA8g61Afa5c31K
I6+XPh3QCO3rTO5t65cJPXKT3IaUH088GEmqUeP+OhepmIBq+pHzdLPebDkL32OQ0yTN3O4ZCznw
xTXJJ+gY4c5HlXWEzPOKoKetq/SseZ5uG/QA3T9Y3hzRO2q2ZUFVy1ZvLIGYppNdVEWpo/lhy0B8
j1PkpLVk2dlJRsObRleBjjLCiwzYNYjDThp0buOA6kAP09CNdBKNdcXg9r+9vh48/M+0OyFk3xnZ
z0egAXGtloRF4Tj6BtttpeZjy4RCVPHl7sa/VcCxi0TMAqASQcv51sTZRhJcgwom71YY0O2j2X5A
jdyVSMuljRCT8RRcvsipzs+s+8LYlLfeuT7oZluqu0iQZ2kmpviGb/Yf2wfJV/pshGJqua8Q0ycM
q1RC0DwsbTIym8VpzOit6E+MQ9DxzOHKMRvPJr7rubpyj1iy/BuDr4OBnwJPrhmpDP/QykX0LLqx
wHO7TuMYiqXiQ+5RkvIrMLPbjfCm+5NyQhF3r1BZvNPW+zkGzaR7H2krf8AQedQiFLEcsSHcfP0I
IrfKESO5sCpsHYPtBUAnkR++D9hbyzF9PDWfSycVFJEP+ehkte0ElamNxMNJhAgCVvPeE5dPEikN
2VGsprBekRd5zEaiN+w2R7B0M2OeELC7J3YnMygNBmCI48KQOOXRI/Uj1oZborg5WuAVII69L5c2
HlmvkmcxWHSTnmH0Y8iLoYSIziOaprHe170QVl+7sKPSuUlv5IujY+9jwd35SrBa2xmtM/SM+srr
LLB5rmryiXGkUOB8d5YLme2Jg6W4zc+Q0RrdjZTLtgNYLjTRu7Y3d1UabyIMlqoBvAc5SHNJ0mmt
7vE6fZNj15nwpRD9xIATCJ5o7WC6URf0TRIlDZ1TzWSmljFaH7hU+t2tpfx4G8u+bQ2Oro4MFOpG
1i2FC/vhp68n9pqrdK817V3/fAuDyDB2tMMMVn87H97OM0TkUY44SNGs8PwRp68nmt4aaVwn2BFe
WpgeW+MglUQVul8oEn/K4nCppEB9RTRL1HlyYQIBRK34G29siIioq03BfWZVELiEXuRIsoU4/Cwe
5rxORkNJ3IjAQbXyne4+nyLaXuhuMPsOMuhI+DYKciFqM3NGPIdZDvqVSr1320MUDnv9vOD37/A3
wiMkwtLLq9rppowkzu3m4VfIhvADuXWO99L4McNSbtg8fJSS7a8SpfATrTUsnBokxv5W4PQQCXCQ
8FLVGTjfkr4iNA6rN6pTe8E/w86wv7aEsVqadtcp7IRAWaqI6JJ1Lw1U/QJXhFF0XLakpkZjhymW
TSFIep/3qJmyuuo5V1JrtET3nC1OPTvgyEk1CoGIRIDd8yX/LqR3MCjIrPeAg/2k0fJ9VQs/3Xat
jSWEV4xe49JAazK3o61V3YOwBJNa2wAuaOO2LynDmZXGysTKssExxHbhAm4wv4KEU/rLn1Th+NrE
QUoRj1I+DJY8u8pkLuCfufCAkoZxaVYE4ZCD/OST+dDW1G8o1f95BuJiMwCVjqM3HCzsHT0oEEMx
MUHeqacvW01HA2iiHGlLt0nd0XwgSC1OTaMaYSnM0yIkOTLoBQed3OG6s4LVVCcv1j0Jxx4KYYbR
8HPH/5cn27BGtFdMHvXssF1EvAd0KuRplS0gDVtkqHKl7o9FPWiaen9DE27V9lmpl9WXBo6MGgCl
OMIYUl1my6YfICdn0OhfjKbmVCXLbCY52PC8BXmiM/6/DGcbCG/QuB9CW1ZaIZHjylJBYHwpMmM9
zQovNXcC9bc9q4vTmXTvxNpygPp8ruQ3IyJZrHpZfgHd3oOFi9Jwrzouc4BEIt/8Ix6LRUtYjMjQ
5VpkiJA7y2sSoVTDQcKCxfOhsiXsDFtzD726FevwgAKK7MLauMXojtiggwPF2am3+1vbcrNjPVq1
GOWgTEL8+J/bdhtoDJiCgJvK6eus2lmck1+bu/oMXqQVkM5CuA7ztHqeYnbAX7sv5UUgx1hv85eT
uln2ZYXQ1zU4V0ZvhAKYDq6yIh6P6OJXOe0hgmRtxMgX7PiywsL4gdt9+vtVZOk8oJejJvzk1sxz
ts5eL6eXLqwcYRjQ2MS75eb0YaRmLd3GXYP/VI7aWLew0k7WkhIu8Kdt3i9elp9Z9z/ou0X4VRp5
hFYGvtXtJsUGi9Xkyk/jI7DD9uulIEgCSLktH5Q8pnCDLxaMcuVcv1qtg/jlcgl6k7LZxyoCWNtD
h0L7VryGG4bgh9DIdxhoXEYM46kdQtdY0BqN7jAdEQ8SkR4aoMQpM2gBt47uVF/5IH09/Gqzhs6Q
fE1bzFmSvd4R27kej//eghVRAy1ot9QUnbVWJkJxbQkb1xRNDFNdXzOQctNYxwfADKEm2CIatxGU
z2ji8Q1GcSOy0u3Ui6ogl0keguGtY8FI0ZPP8UKijTxjidTbubV1UpOG1oLEjpYrYDrwrArV5O3H
RnJxoEfAFlKdc5AtkMclKFZFGlZySngdv3hAJsMQkC4fS1XHXoWr4y7mz/e9fiTgoAVUVz6eNqfn
tti4C1Wp0X6GNlCgbuTCKd95R6FU+KhVUj2vsYv3psN9uWyGEAZtEuTIN2oZEkBgMiWkHYNUx7ur
Ls8j46pVvCemsRDRnRgMCGoj4AYRMixYTuXfKr/3OafXBOSOVpcME59NzIdVZLzVqdMO9kM0MpyQ
SJw6/NTCtoxEaR2wIi2SjNyOqafz5KXdzFxkdQxTBFihWpqpPzp1d6sPzPEDB96q89zF/v15fDa4
GXpSBYv5lJ7e2Htc9FaNeYelEr4YOYbgkqPqkeeXNJ9AU+8/lct/0q+Pcj6bcBtC0aGnVL+xKGLb
zpRobuCJo3m+TRhL1qjkK94Dv0p0XZUy9zpVmIKTLJFfIhf9NUVK24E/4eLKuOpNspZuzh5I2yMG
ySFeWwQf7+cpUJByyQ6wBR0Us0Juwqv+UdZh86RjJPLnlpnpILaAPbgligtbxXQSHJi1hIEIjIJc
XfvI36mRWbHkG+fMh+vtKvLB6VYcMtzbnp7kWb7Gjo5xVEOWGT1BaArwhj+OFmDFGf+TV6N76qjo
SAaefQ882Wpz6VTAsGX+5G1CFHx4Hyq4+nuBWiWcDSdFFpfJ5zwd307okCEArfP/yjXFKuBqmO+d
5h885z3EXNHVU0N/uOjPWQCvELW2vHWdnTF7YK8nyuLZ0ibbEv9u1kgPw/PpwlmEa0wobNSfA/U9
IReC6WvOax+1vDLQH4/E8G8tBIhovv/jkg2Apem9L9ROsMcKDAr0o0I+kF6RhFJ/r2CIJI+uqz0J
ATQd7tRQnpttYmO1vMazxx1JJjz9SU5mQz35HwQ5ur31xMMXCPZiAUl6jcgQlv4EJaM0I779vA5e
L+egtb7R5fXAZ7VZZCZZBESpfXTGfdkK577ouEw4Ea2Zwla3urja94zjsieZtzcAwcjSI02Fr5Wr
Kau4DSOM0G9Fl3l+Vb9J3BBZ1nkTlSelbFfPPRvxkr0g7WZ7PGmEiP8J0Emth93MKowKtZVU1O/u
6h54H+Ux/NbBH6CuAlmeeC18eSE54vVD7HdL6cFBbhiUtBfolzZmMeMp43CRqNk8LKHOfg9N5LFA
yEEW4H+PRxvOqWECJEHQgssgSnqghn36UVTUMKEM8TgwfX3qdWaKqz32xwuZenmvZgZaXJqU3ddW
dqw256j361p3UodW3S2FAmfwg18nHym2vhdBIaDwUomWJlm7yPPVxpId9/H2AJq1JOmOtbOh1CaO
DS+WWZ5ZWyJVjEKisLA9QdKfzjAwywfkI5AuRKKPUc9dlzG4YVELC2kCtfHL8ZXbmyZHzmvKhDMZ
Ect1UafBSpf+tw1xjS9HRNgvWtqHRCYOXvQbJCUJqeJ7CqgrFidy0UE6E3ol8cGS5K+lYGP4bzTA
dp2M3QtOLjnScTPT8OLnPtvOrDNmSWqACd5RhGE+CmwZYzJrKqENXI0mLT/L1/MvyRQRG2zcgsWY
yogWeXEnqJtLM1lfAEMVEqW852h4ostY2IHKZsOAml7jA3K22t1USDVoVI8Cl9Sep8nPEJZB67Dj
ocPF3sZdSL+dW7qLmuaSQxNjnoLBD3krzztZWf5zAQqG/IYR/CJuVr3C6f0CqOwYZUqVLzVWgO9O
tmcpWnTD3bnMbKE3gb2UN1JiGd+P+Wk8CgmB5/DSkDl7Uuhbgd2u/pBdyBe1CrTqmKfI7Pj0ICs6
vYhCxuTfrkTPUU6zXdPJdm9BPqy+rCZnoWddl6yibluDw5QwaAvb99lbbfAsss7RXZtpfe5YLmgw
BvBLtQMw1FQm4El9T/84N4HjVO/EIb5HFoLyurL1MAp54mphJtKyDr2S45ztI/fxHr6z+ZdElr/v
qCnEUKrSEUmjFr+8Mbyp4usd55aPILX36Vlx+VYyJLHNSTtvxrtVoZsoNAammG4Dtpj6O7pgOiQn
IGRZXw4uXj7Qz1gcwGBJsfQsi9HF8SV8wBygKQtoQRrqGhRDMGv3A1cu0OQB7vbUQeaMIxfSOIpG
EM+JHuRPj4sW0QbAuJzDCXSe1zD/IY4JO9GZ3ILw/3F5pjBNbHp3ml9JfnzJuN2H7R0uXsf0cePw
OK5PkVcIZ1fekeSudgfACIOSw/vrhwWk7lsMa96iaALFTSCtAJII4zKIJveNfRuLLB77h4hrgs4L
z6FLw1ymDhDyBjHRSVjPQrHNix0C9Jf7sbO29sN3udYUuIeaJCsEw3WOdiZssjpgNT9/RppF5qew
32rXWg8J6j1JhWQt9ECgoE2VHJnUe4hWKIvSY0WiXAyw8TL2ltjwk5P8fLkaVjDap1npN+18Ix5D
VTNp6DTkxMWE264IlrhUQoCZvZMCaZN7c+8rkb05eSSqF7a3jMFpCs3qltA5BQonFPbyahZ7WM3Q
3n9AqdiPhFDPlVoPEpXZn4qzRFdxkpN+ZYHhDa7yeuL92WB3tqXt4oOipErjGjnFWlLvEIHimHaY
7m7IFm/I7PZpacSNM+54hQHwok7uVe82PVPgHnP8Y8CyKUgGfMUy7EU0i0PDEzrSIEQD5cjabMUa
JCGmML5X3C9GPQ9h3uQROPb1/NjmIK3c0rzddc/73Ef5zME2ONSGsXK2RFt+1x5nizh0DpTI4IxY
PpQBhcqj8oGPjRhemX6scPcDkMVlmiRWUJywd6v5dI8hEDCS1TCU2Xp5W3NbHtpxo9cZtP8C0npB
4xs/0iyFL/uWbxeuT+a0N4eitBfD2ctQQ6NyBUs7SwsFF00zob7a8Im4Gv0m9fSqfCw+fh5/uTVa
jvm2/r+ktA1e7Yi1nh8kRyEH4980zStcSmUQWoHGtJA8vV2SHtdn78N+oVGO5aftuMi9LSQmQ2gx
DzxJQBSXRk9SSCCCldszsRVdgac95J/IsAGL49AJIdb4NvVDDEDBslhIyoOkcNChMjweGO89o1aN
nqbd2a5tmYgTKVm44WF1yza54K3rlVywqDXUrBGSZrs5SeD8Nf0tnqrdzQu129UVZoy1unfrn+j+
EK7fcwSZl/XMINfeBsynLzLnhtFFCdRU7Ch4lEK22rxKf1lYhTRo0++BK43X1TlmjFebzQMLWt72
4uyWk/qmgnBgcOpVfSrg+4cVG7ECmz5LJ1ynl1Bt+85lnLn7e+GsisiiyyrfsQo/p4yQ6fO7TxoI
LpvSnYrziX0JWtvI7ihqE01Xn+zTVpUAINENk9XR+TsBLkvQyN2edmwpo1AHkE4cVnqCD0m3SV4O
XVTD8uDU65cStbgosfuwtXmBUPrNKwfvzzA7CXkzUnFBdIiRn3TgJ7G+Ggj1kBtZLqt3tqdjURfF
AZQtfGPphVaTr/eDbC0IQhzYMavj1ng8+3ERHOBYqNVmr19r0vMp2BtPgKlrWvhHmkjhK6SWU4gO
WOoZXa9Bwx2e/KphXfuxrBnHrwFFeJh6QthrrltG//cKrJZrXd+GMRsP2l1cv0FZMW3UlkYbmP6p
0VcpOpD4Opq5hL+vSpAGhCs4tW7A6IuL7tuNEXl8axmjJOdjuFy/erKVMu5p/+rXjMCmZDevuf1w
rTECPrM/2+7kMJgpobosFMKzG1/4JV89LB5+ei97JcCIvyWw03bVCdbJ6TnmtJPV+NkV9Hmn9+Vb
ZNbl/MvW2GA9foCm5XVObZic2jAYr0GJY0XqhCdHHfAkRrkdeCp+nO1zAuBOHYe9NhzAhHaWj3oy
e1OZnCTBCUCvUZjvwbsJC8ZO0ypoWnQJLqMN+ZmLhWoU3IXNh8RRpXM85uyosQC2zWQ6WgfTOCWA
WsCasg80TGAEt86ciN7S8IwE9cu7cwBXBBcF/UL802yvin6BFrd8C0iyfdmEIJu2EAiX0o8M/FGG
iMeWvp77ttMAvz7iJLZU/yNCPklWHZXvle1raZrDGviKHlF+Pmg8wSzy5iBvFtkg+OKSYmFExA5L
7Afsj3JtliqAdE1XtEWPtDiX/wsO86jnVh4wj3DU1ec1lxuUPTkqHEXj3DBNmBEzMM1ti2KlAETe
FiQJuKOjnWaXXTzccNlmz/egxvmBNuDtOR7zKimEwCfQBWozrdtS0eDNVfWxIZRhTmO+18dPBexT
4jMkZi3Bz16vYu+wpE5WB+fxQjgElIO/baEJUBCw41rocIkN/sVe97KB5AeqI8sAB8e9l8lou6gs
qEOx1BMwkP5vkWtrf3CuZyjLVIiN3VI/eIu/UeL0UG+Wogt89af+GQN3YUSRRW7+5sVAcbRUj2gp
bBHYE+s/5RzeB819yB7Db503ECa+EA5YZclcxQkaDKoTSV2A0Lp99RFE9CZufT+ZE4LDEPefzR/K
BjCVf5N0SMWf0Jw+Ys7HNydbtfLBaaLSPXl1CA+YalMsj1sik8dxv7YRdoW/D/UEdLA49nV/SkJC
nBxpk9r0kkc9yQcxdN5bhk3Leau01YCONNHe7Y75FPa6xqc/Gr7YejfFZeFl7FlJ4lpa18Qzo/CL
PxtyHl3XPjuW5E7URxL9b3rqv3b9ity0e7pvPVaoTfiPcvMSHIxswWKLi/EGD+RB188ILLPYAR05
o9xjXP2qGg3uVuc1Nx67jn6MCJHCq3DkPCNfQwzBvBKIGUbExb3QD3uF7Icou/lB7M5MEDnlHT6j
H0bBDEPAo/+faWkBE0mYLQebabNzL8gs2yA+32LRCOtlfW6j8XdV/P6B2uhdwbbRuYRQ2Uhj1Cc8
90CHQK3WNSL0yii3MUOhXW1hw6wwn+0vw15/GGBgUMJtaOPVzx+9XoaTNxIpjsD388HvfNvCbYAt
OY4uT56QrNEeVjEHErER09rXk6JCeS3LM66PyM24LL5W4zYTagjOaQ5gQwRtXgvEaq5R+4eSXylm
+JHC6oC/rCZHNymRpxB8MyM09qDGfph8IRqeITvI6esL4/kQgTDEoREb4GKg8n7+1skqcPZPvPU+
ZzOh5Tx47vc9e+OYguUx40ACMmBL6NLgV8AOzsyOP+vBCKM3eH+aDoHkCoCwVCmIh7KVc/ZeiGOd
UbJq9UWno28Sv49PLq8LL5uRqZU5jf4DVjRkdCG9LzHYFYkQYHoPtfN6Q2l0HI9G3/pgqZs4FFe2
Yo+D4LwyMRKTfLMddWlWcDilzVQM58C4o1Vs8l3kW2FqC29UsdR3faByHtLy834jx1Qm4dU3fI9+
Qwpsz0gHvOnY3oO48mVYBKTo4ble8C5eHWTp60OGOvqhxtJ/SbuwwC4oyid5mrGxE/tx2oZy4QcN
WeCrJqOP8/CxKjVuf2PzXhNo7zS+ufE6UlP9tGiDmsvaPfhdljYF7z/OnVRkmEla5ZXx2Pv8LOxl
Gyi3IvVlF79nMr7WGzNT4HjOrFlqppaB/LO/3DzWRrHMRcn4owTobXTtTAWSCNLP9lbJw/7/L0tT
+iVd4a8mNCR0E64SQyvGjtYND5MHam5hi0c++aegTaVfjPWnoEO/IYZZpy9D86sigEH5wdhKC+vy
YXRHygSiMzZiMTdYyBm35M1oa3CUZ4zPFHqYIUwKM+NgVLZrC/cxJmgEz/mrD0rjQpUPKrSKbWat
IjROCZJjyv9F/tr1oLjBZDGFwbMoiFNFA3SjM84p33CXPjmwpPHOTduX41KoeTVs62ZYcJb+Ha2f
PZPw3DI+ePxWb/ng+27ulTvn+xwgmd1aN+3JNEvAMchAlHzje9MKZXTi9C0Zr0Joh77LeAuWP6RY
pJYQvCKQre3g4OmcrQUm3KNlbtnwnIgaQACbThr0VI6ELbfBGD7/DT64QzhroEfHqIFTsri46L4U
7NGlBRG+5L7oXblc5Ja0J8+jzItnq6jOSW7CWY2mMCodj7eYqrmnlIrmPrOIP8xZ/t7whrf5yaJw
X8pHWmJ5COPE2VrapVbAIlRdzCObj/TlSLCj+xd2eBv/C4aao0fpl4HevgUgIq8VpEZyM5JiKgbi
ci/khrB+5bG3SYOcjb1fbVTJoM8NEh0r6GMuFHBIdmOfliRmKtkum4f4SgbW5UxyGUQKHRDSD2gK
hwYoLxLuaon5ytSvwe3YzxjGmTDCMts/AQaV0WOW17alLMcDMACTY0rzd2GMHD2M0czeyXS2ycND
83qqINZo7nDTNHc8WMZgIQcbYfWJDs0Z+NuPbTeSrvslW0eX6UHqevv3Y/aPlh76TIwOIhoz4gLQ
ZVV+cbchDHCdcp61f+qvVCo5Na17wSKgB6oLKIn/QviCQYhUE3PFbfx6kvIX42rRYiAJxrp+1kWp
2EJ5K7nIUdLeHjyZrPeUOXID3B8F5VlKNZJzV9NNMxdFxS3mg5MmL6cgk2VYEzkK2oaW7+j2e3FH
S+dUFmWBEi1ZKs1GN5FbaTFHdPjuXc4hpP76xpfRIxynK9GzoEvyZg1q7QqTn1UALjf6aNMZRB/c
PVIMeHnMOzDn2l1W4BTBzCcgmzgr0a0add2cjIvCh8dWaGzvxiSD9UdUQ3AXK+oKOIoz+UXJJIgr
9ALc9wU1qvUu/8PSkOoPtH0bcxvLViCXCmB21EFm80EQ2/aFKpKfSgbVpwP0WghgEqU15FHO6+0Z
MYBWdNmu6BHIqJgD21gnbZMs/rTsrD+McN2f4mq15a7ZqkXk/rvXMJiYEWxjxmFxgF0wml4vTrHz
BOER3c4TN9jtcsZQFF2ty2JQxf02X1ze5+2Xx9mczBG+YEPpapwp8DwjDLMw8ETpnpiDCZolqdVU
NHwDHtylVkwEb+JPQf7x54kulbtlyjMqQvcNv+nmpdgGu/wZKN5tOFlTECpm2a8Xguy/ZS1ZcvDY
6tADZoj/f8/dXKJjCAm+OV6vjVbUP3pXaV/LE/71uxAeL2353Bs9XjicDwypf3snDXpCYBU5/hCg
NrKibj8+OeJmX/50Kz9sPS8cXmUvdxYXFRrMbUIj5AVFX1QxpajlK9PSP6eSbozNZ1hYnI/2s3F7
iRa+laymsPth07o/aSaT/vXzPg2iBG1h55vt5mBlXQkfwN6CB091/xTi7HhCx6ooAchONrs+j+yV
bwro/OQkngU6c2iCZR2S1PoSRKmwkKgxeS09T4Rq90RM6oz225TJziZ4cacjembw3mrZrs4Cl/fR
GWGUcaCBV7/kQiq8OKO/2JKUXPGs3pb8K6yb12iM+IZmX7TDRYRf+lAS3+N+3hOlL4kzEsb7yY9+
qk1uGjrYkPjsWmUqr1KYgnErB6vWLTy8EN8N5GZGJu9S5oFKLCNyEslxlGMe0oTpbdtd3lII3d0z
OYdEqi8n78Ox/O7AIkrjRPnG9Proc7lPRNfNR6lJk/pVWpaRJ6QOtj7oqx3TbYgwovnjgQYtQnRg
nyAtWJCzHHgHJ5OvFf/rdWmx4Y6sTQPYJlOtAZvwlkrcvZ2JzCanT/M7a0un6oOmEaJ9S5vJMJiw
vmQceN4NP+qFdAaG/Ulhg5sNvXYveq2Ijb/TrvQ+FlnlCqaIp194ajY/tkyZrM7Z/hNAZTtSvQ9z
I+xK0XRgzc6SqlgjnyKSAmm31DwLd4PAPspMCvRyXyaJRodPzICcIyD7rdl/RHrpMY6HAqtzUCAR
vegMVpdyez1a0rG612r5PrMRjoG6p1VAAAxldiCe+10FghSXeypgdaDD+EszZPQqSLI+g8dfxnWf
QK7QDKEJt8Rdj4cGhC15uUwNqitjZ9GQFkfDyfpJGdrINvNdBBWsx9xjl6R8mlivtS8HSonIDDpM
05dajQ/DSnrup1CcNAYuAxo+sMgozQkJ8CBN8HN99/ta28heCIaisSjYVY7P9CSRHTdsDGIuKN/m
7WQq/Ksry38opO89954oIX56iE0B1S9OwR1VEZhk6nJKvx8yzEekA29G+nMsMQrPy6TeAQHb40Ar
hjDU0O65pemueLniVP2YcR30Q5d1LvQeK4jMu9IAMquPUPvpunCBMvnIn+Fj11GMrZAl8Yzoqc1y
QqbuusRpBbN4sq1tZoBmrLV2ImHA34DPx1kEfAthZ7gYEfdicictMqbb5u/pm9CtfyHWA8LZj4LD
nhOxVhppPt32G14Hgfczz0AGqLtVWsXXv2eoNiki+a1zgptkkrdqOtC4Ju1BQIWiEHSGyG8AXHLR
ksIuI8ntg36/TNrKAr4N+vReNEzQfq46+HpWfgWWbCMdNFOkCuK8wKs7uXHgX9NeW2yQs7nFKMDp
fsGCKwLSyaUCupPPfhkyTS0aFyz8I6i6r+eBeHo38go9n4nV02ivUJO4hZFJAgWNfQYZC3w3snyU
WPJ0J3MYZ2wQhKrWuPjaquQOUvg/TnSNnysNbmxfH/DptHyuY+h+wMRDfw+RjKrtTY4/a8HK0Te6
ffQp5jzeRJAiYkJSirJo14QAcYkC6moPzweELC/1LYrtUtwBC1uJXgMVG0cCqd8KyTD+P04qrqLg
wQrtXggJz2IDK0s7IBRsOgV9HFK1ilrPnQI8xaslNRQMn8+6Raz8WUCuZmITsngqA9IEezOU1C/b
FviCxNdA9U2KnBy378nf568Ks51enGSANdj3Ze4I+VX5pb/OIa6NTNIwRjVGqBY7rI6B7OkyzVpS
BoURq5qtyPSPXlYi0cfKqkWUm1P61sOzQkANZRnbIalMV2tmBmVMzZ+rIoJMlXQM74yYl22xZwen
PImJGAYsNxRlu8fRrGxGCzKhDnHXD5pQWJd0HkWrG/8ouAZ7YHoWTjsjzUKi18D32jpoNNHIdUwQ
HpD0VDVLkT32BpSX4sJDeyFALPGV+g5wntYofwkBjlppaE4fmxpqpFvyM5YM+8V22HBr9fZ/QzK0
MHq0GDdvrb0Qa98j9ZuDWAEOUowdX4GG6OGlWiRrRAQ+xNtFmS551I/DrfpvrL2SjjLgNHLjh26x
pRlJZ1r9ojp8bo7QGcIAtdcM+cwJMIuBR6Hvcvugp26tKMOg9tBZPalp9Hmm4OSgowYN3okPJlSI
v3OP6eWB+6ndgVezEmP9HYxHL8RW5QsQT5675d/HZ51aU11cyCzXlGMK7CZW9nUhWBVH3mcMovSz
dohb703yx79wkXVtjWNZow3pnwt1LSM3h2lUTXRgQqMwLuQqp3HJ0bUAPh6lkuJEqafuvXs4JI2s
Q0nCAzXgvdVZeKOiHxNwAcfeCurXmQSaiwN+wrhcj8VYphqLMAOMBShIXvv/ANDYk4g5RuOdLa8j
EYGW1b/ufVSA82rlS6v88MEbWctliS5Bnv5mVPDDZ39YdrcfFVKLweaPlBL8y2zEeYpcSrukzQx0
tmtl6GTmjD5HeCK+rwUIYk3iXRzq0gPGk1snWOiRAMjRmuXT3R2R9ooMnIpVJEwTiIy3752lzIzY
p3ja0w6EndBaWeoBLEyMc5HHlhPNtRWTU44mwWROOJxSWhW9GD7lB4KwIUlj/tQKCe2i/mxt2/PL
vb4SbUoKs8HsK+D7LVr+BSUez+MAAQLQNRfmD7LX/Bnvld6KHvqkwL02+8peMnMxeInbo4REmLpZ
VFJ62vD+XbpHQx9QsNcNVKsnt3c0p05jmc/zvfQyxzCTMTee9UTXMx8UUAjBHMcC1Gn+QwrEkYvQ
3Ag6Su6jFm8jufIDQdgNBO2caf0WaoCsTxZYhnlaN8AQTs1hWWSZ7xPi2TpW46m9UyYhywBtmrVg
IaRVBhd30a7YKPepQTStqV0SDHGvAP5kTPjfpFvzi4BqJXMPSUVb2gg/8Mk1PRvQtxZCoJDzkY9X
/r0a3Dy9gKOtwGRlbcm6ypiYyfOFImxfuxviIaX3Mt3cfuQYxXU1zwYWrzmB02IdVs75C9uYPNI/
KmDMYOp2tUl2bJ5GA5KtJbmtz9ob4P1pij63ciECTZcmq+JSzk0MZNHkXTvv7g/4e7/lUyAr0cjd
7fa4pbIJeaOp/iTez4ji/OWvfCYldx+7ijU0ZEumo09risJtF7F8Cf9YeXor0QOPVpBIM6dFUPBW
GN1CkyXqVA0J8sIRPSnmbpO9THPZuYYPWPfk+/0d1nUp0o3/gRrTNXLidgClvRhdAaYKxAZtjFwa
kvYWEtOMb/ekZVEjcECpYKHJgHOCtNlQpo/mbpWxk/MaPirTP34k2A6vQ9hZo1bUf7aJXt37AnF0
+BC7VVNgPq6U9sm/rrTvCfhfrUlxnqRt77ZtWPUm6yQ96Whtr/RnOReBM/tbxYuTUO1aRMHGJC3H
zPajFWdiAtC5ogSqyToW3xdhn/sh8Men6I3pYQ59gzz5Phun8drzPqlXiwWuqPf9sC3xu8J3R4rU
yw2gEzisybPYLDRJApE1Whh06Nr2gwP0Y1D7YoR3csAThavG4Apj03Xs3GHyB8fRzZwy9r1lBZsU
DxYqNNllqGN49AdqmKsLtyRua2pcIHydtrE2DV+1zJUHFeJFW1eKMzrYSAjmwFw9gTMDwNHx40lt
Vh4+yPWgueGoMjAgvTwUfp452/nV7g2r9QMKUHH6ymYZEh9zzgBoWMIenN6DM/uDZn7haVyJaJi5
w8teGCPL6mvQutBIkJU3H7V38va1LgGP3gqqhVwCs4oW727vWe0ez31R/aBCRX21VE+bovl2vPJl
BnWVI1wNE1b8HP4T0pxBRhHcZgR04gbOg/rMl5wAb4e3jPwYznXLBTLfI5kPLKEeTASq7XfFcTC6
T9IJz2ucvlZpSTtyTPxClKSEJsuKbjZUHsZ+MiadOgZWOwc7+LIv2EP55ji6tdXQcjOqdMSkq9vq
BQkVh/SDnovdzaA4kO9NQxMkafyEN5U7H7fODpga+F06NgQIhTl97elMNKuFnTm5joZeei6xYcaD
I6gsb4sFvL+oYKqM5xAOQQAEwGNaaE/4MBZITr/JAvrPIXQF9SYlmvuqK1v1IXz9X3bZVuo03+X9
wDBrg1WlAm+vf80255hs8502uWfVnYYecDkQpSRjJ5YxdEzMRwwtlkpZQIjqWGoFtjJMlR6H2mQ3
SgyhDq2Rc7NXta1duafaiOZyV3ftkBtzYrNqT0LDHkMvMhgALlUbIK7TCtokGvgywibT+VvLSayn
yPkxfCa6//OdEwANayh9VVVyICR/N/wt1tu82gcON/bYCPwBIg1OPN2qFnIEsV5CQPFwpf0fYOZW
Yio7xbCo3MLpORfMNexQywuQgteau4ZCMlvATNUyccyY4uqymOav+O6YicD8QZVFoCO1k3ocHF+q
fGBXtIhFAZBglAYM1ue8oXUnXmYeFQh0jWIGTemxM31b1hsOw4JRKDvHZcf0bJ32boDSgxuSHdjZ
T1Kw/i/t3lPGWBXtYbPo/96RfFcsoJC8WBbHqbLLU84eOwaS2w3+NWFnu1D89It9WNmwb0rUAjye
Szwdm+LSRS9f/Kb5RZYKeO3jAdy96SXbcRUiOClwgVmDwljpuwE0IA1Cdr592L9rhf/dBOHeUSqP
PWqzz/z4BNk4AVC4kQ7OtakVIxn5txoPcJ4Lm3cFl6oAJ25XW/MNotWsYFwSUehk5Zu7pGV+Xaqo
Pol4AGAOpTNEt0P6MgkU09fZZATvymCLkOQj2LTvMCblt+kMgpn7HNFGW57Noh8lNsrxxX19TDqL
RoYGTQA4L1uHRVk7ugQad2RaYdvFscVJLalijkmih6nlKh9CddnXwL/717dESjsyeL/WNC9l/dli
1D3qCCo107WEIGcSWpKoRxwMSLDmKfWm1gttdFeij7R49UyZl0L+HhGSRHe5gyoF0jRi2mekogzI
K7zzCDJoMkI6QyzbvbW07vkOAEEuYsgmrkr50HARmp4j0x0zA4TySDKkVlpkA5PiIhpXiAz7P9+a
63vv0EWYypHJqYJvLdfIYNI9CcIegwjvgW5IbOWpdF3D6+5bd1xoRl9ayF+Zg7ExByUFq23s3WkN
y7kMtT8NBvdz830YHNBGOx/qLTheAmLqbONd5MiN+PkCEfePMnom+PoIgj6B/9/kcn+CoMIbYB31
A/bpr4SPPdY+oln33jH2Cdb93rvd2m1uvSl9VskD0abBA5t0zuG9/xC8fqGzJpaFXoZg3KRuyKZC
FmNtZxcMEj+GSzhPeHV6vh/kMBk6J4rvAfGFueM8Mn3wNHaOW9wDJhqE2aYdxZBbSSu9ebWuwgDg
PdQTtyyYic4bX4jj/Jsn1kmDXnYzr52fGDNqaDN4YW1gRpRSu0ckLPP16uvjbfaZfdtM8cuDMAYD
XBhyaZHmP/AqNrYlVtmRBF5/mA0G7aaOS7iGnsLQmVuY7NYIJZAQIE9/zE4fIKErudaYB/WhyPJ+
6sSxO+Mt/UDWm3TBC5+9FB1Brt97Bcs640f4oU5HIkP4Susoy9rZY2apmjDzQ/a6YeAPR8HhvoMa
SvktCs2qez9oHbTQ8xxBm1ict/1fhkoNS0uxq0ti9+ICcjBr6Ycmhb0E+TznmxCD+XxxcgPlCIlI
wNAXENxUqodeKQTGAno7hA3eu3QucAC95dknN3uJgYYq2Sh330H2UZOqswLGGqCvzC303xK1k5ev
H8z6IrtKNKFLS+VQn2GnNy7rABZ/nsY8VaqsaKmFS1gntdYZCxzquPinT9JHqTUKOuRUwte+M+n/
bp/FjvSxGJAOTi4J7pr12TETOqcIKLXggyBUm07RN2ZTZOLoRpM7gYSI6sNm8QDFGI0+ObRkw6nr
+xWTUps76rKQwq4wLbqyw5TsgBqVwy2YKclsUecHUxfIRas7robScYqMUTpP7tda3my2Zy0033wg
jxrq9OSHT1fAdoJ132NEEYViQ+6g13uHAGmoI/uKaZ1nj7DS8uWw4x9r9+4L7Z8PI4WZVeB2Yww1
gs0onSNcHuEvwgwFAsIBsunpRJNabiItdQLZIL6PIM87tMk/C3glt3jdpMXmd8FZkoJqXtAGyN/Y
2pss1nSjYEuKG0tAuGY+xIRonbMnRqJ9ClEKh3df8imqMqhnHeWINPxUQ/u/YTaYyERqwhkD5+db
6eDStbZwbbFeTjQxUmABHw7PwfSClPv4dgz/4498/+L4ro9FcU1xYFfRqwgGh+9Pe8rt1fzQ4btX
hDGyhZZs026nWCzJqjUTlmDYqvCoZsyZ459OR3aeQKq/8Orhvwj0QblF4kjfkLtmUXgTg7KK08Ks
khxRnJjG+wHPuD6mZN1edpYUC08uVXUz5AQHhKUsnBJVNZR6tYiiQ8mHY6NAAf4z9t82Ezra66/j
YoT4OOBlfJbrfoAyI0ZljKjutwswn4oDXanCbi7X8OwkL8Ki0QnEqQA0oBTyKVtV+oMMtZXl9eIZ
pef+SDhp6qQUDzew77IEQM6ep6W5uo5N6z9NHoI9PUJkAcWVyHGMTs2FtWlpFP+mLFmmymDn3uH+
eFFFLXa1oRC5feQZmGB3h0k4R7JOOpFtVR0RVwMxRiEzTN5G4lYK4h7jKdMlxedr+s4QELfme5X1
CYdHYHM3tx0aiopAetr18xOFY4FQpmdNM/iV2RAAQPCPDA8io9wFZVs/xethYTbfs362VmhOCRL3
yfELAmfe+62BkfZGyZ5Wf/0unAsYtDT4Q5X6kY+LupVXqkc8OOeY9S1VMI8NSH8o1/6DYA10frED
LKSUCp5Fkh9POwagjOI3GnKZ3LfZ0g8ueYkjNGcDKLRFSAgC8Z52la3l7uFX6vbSTyqy6XmHrusB
dCCuXoilYLwdtjDFRslJvvk8/DIS6McujXgis+yZkiahPoBpxEe0HbIfeWACCH+HQ+OO606cIwUs
84FHCdSgWgSSmDAi1d/+ufadM3gxX9BMtAQVoeV+TFEh5/VBih0L7F94/y41jlkI63BKaLujwqHD
DXmtbpFSruay1PDnH8ErEA8RJLsjAkh49F1a9drYFMBw/6i275ch9x0U/6EM+A//KaVbHjncDyOl
ZT38EFRi8XcY2wt4nPDU7nLZEWC3gykgQOlzFL31+D1LlBRDyQq/fv8CWPoIc3Fay9zVeOzZ7aT6
HdouYTXIjcg4HPz0hAMaMvC2q9xiS3EAscwR2dOd0I5jGC7baLzocMmwDX7+Uev8vc1GS34RV1SY
FtZy0iB5uHIOCdd8rxbRiWsrVZ6gAKIdLcwVcxdyUwjyR7fekjVW6aD2c3ze2LspLNuP50tG7bF4
OmLYgewAQghREUBF4Tm5BLtejOJ6BNttjsHSQWueZ7WZYr5Bhm0fT5XsZuPeYL9ZtyLJaiSoGxE5
hmoFDvJr3dtMzPd7jKSWoqClwzjh4brHqFnWvS6txeE3OQhaj8W5X7ZHWB6psN3UNBHGGxYNEaoY
g+Fuw9gDVAtWEKFW86Js2uwtoYnNVKuCdcRvQdMwA/BWTu/zIbcRgm7nJN1s+UIyjPCGefe1zECL
tKcGbs8gMwdVtJMqJEMXu+XpMdk02XiQsjAJWDDtIU+SC2oAlNC12AGA8j9QTx6Brh59T0spGVke
m8uHd7C5bw6WNxpm/TVIoB07aSJUTA7byp2a30UNoTSgL9dMUckUPGaBUt28Kp5nvWmJdGhH9mys
ADD6XyNvS5BSrVGOYPrzJH3fgcVs8VdZhYO8D+auSjXVFSEYpYhYRv05sYWDvnIq0vyeNwgaE/Jc
c/q6sqsEdlgm7wO095KB0z/9hAEwtL/PGRs+JjGwpxtizdjd+r2mNQOVl40eRwIu6K5RxobJVXYW
V0TBvV4wl56UiHMjkw/i+ICKR4nHswGBDGdyvPcua8oZWfQA+aGo5WIs3Lc1RWM28kEXomJwN8ft
FmIlWx0u7F8qQXPoBwgEaHftSaYNEBEA+tywNstff6jWiHNt5I54YvdUDk16JSNSI3BgZV4HrgEb
USTq0rbr4QscyJacizgHkk2wRLpsBqxSVhUSyta4ZEXrh81Y8PWkJRQDor0sci/FWpbDHHXzYwuD
DtM1g+s9KVgghgKzaA3sGuBwIwIr2uqvY/FTMXuIQlIeyCzfIwyh7uDdWzNKaHruCJ1ryoib9oii
U3EuqGQ+v3ZpE4wMZeOpYSFXFIVzlQ19AqlauZ0sGiXKv8E/syJa49RfenZuicrPpc+wIi4Ne4H8
S5ASPd7x1g6hQSU8T++49x3k/3wYy21TXim+7bSjvgE9RebaEqjulx473/nV+iXgOQX55X1/pG5z
Y8Sr5lU9AOvqs9uOvv32LXxi/XwJDeSlSi7IefThyn4tKNu8VPLOKpS4zMAXSE/SMs3ryHMnoF8I
6sa5UGqTx9msBs8PFWq1ux0qt9JMqWIULS7CceHmF51Tyz2lVNgtuui0ZCfbNKybHsDwMiDXViVN
UBJ0zkZJSS5y5dKkxcBnNXcYABI+1/pV+lPQb7EDR6z2PKDEX5PQof/0Re+LWkaY3WuTFgSSnjsb
zjTm6e49XRuhNhwQSX3OTOYtbiDbbxlauLU6QUCtESiqiwpUL0iuSgvvbLOqD2MEnS1r3zTGMswD
d40AbGmQlL7eQ+VMw3e/l+PXEy7NG6GFo+ZvAud2m6KPnUHXg3jansh6SACx0JwTpgtVqd2dQHP6
WyXMmgGg3JyLBdvX8nW5pzrYi2aKF9JZL9S5L1Fn2ryyyw6ek1mf98u9c8FKawKZhfZ0AASlTXbP
sog8wB/Zxk18GnUZjpSlQcCN85TYOyAfKOo+PpB/YBtBYUh4B0TbZn9rw9MeV33bMw+FxdEyUi+F
OapyiauT/mDVvFXJBHm1sG0zUyC2JFDEMfA3Jzob7o+o4Td30AZJ/XLJ6n+VUxyD4SxpBiLshuVr
zOYL6g/xNsiljfhdSuebI4LyNMlSQQd0h9Ltr24orG3zZxHxIPDxPBYzvur6Me7hnKzha11HAgk6
kJI/Z/fWbQZhcTqm2NuWnrlpMGlZeM+M8r3eS8tvXe1a0ggPJaHpM20bMZUFbdNCtNaRWTOVeN2s
cQm3jR27x/1Wzt7XrNgDOc0vBGDPcDbQiF+Kv988gfsXtQRQyU1KJklgtouGJfKsYLPF50UVtr6z
d2ZXlpRh9iZD9ixhJXkwMwzk85qPuDO8k5HRcEesKsCef50oPPejEJvBq54EUC9YwttubLoJcc7N
gIIaH26KhhWo9agVrZiZ2huRntxuM/Zu/+vgqTsn8IqzAgp2p0ZuQakxh2z5KqHz4V9VLqDOmBU3
fHpDTDTAxzwx5OMWZOUcMnQV9FmiAqG7YYdJwycDoAL6YJX+LR64QXozsm1GSeVBahnPqZpPTOMo
aLoG0fem8w4vuPk4GNk/73fClaZF6o8+Woi3wuaXQa3XoXkhCKLSvnSaxkitTRMHt39PTTQ+zepx
ZZo38aECXJcFzV3OZmRY2FHG8gj61ZrR0pV3Udtr6GJfznR0+EIdK5mAJ4xJZ2fMj4om3RGG6l/E
N/8MOPgedSg/QBZG+CTx/34Up1uX0WoKinVaoIbcnUEYl1yKAnAGL4pAbhPAtTfDWe9pjVRpYx6h
mq605glms4SjOD8Dv2X7Wga+tB2majxq+i+qGRr6roHQNHkjhshUTfPmolSaR3eg1eAsEkqsNJFG
xdKCTAqFvv0X7HTC9aKaBDeneFiRLypTtnBSbrT/+Oop+oTCBpWJ6ZNBAoYdJOsISGf2gyCmNNl+
q5zemtegizho5SqdsGk1O2jWLxRvqeR4lmw55fofp5gpToxuUAFZXnEo5blKD8ikgO7Zvew19iuA
mMlpG9AM6WaICd0cQbFLisYuqpVonYLuuLnCJvQOBNNnf9f/f6bwGkUioy2f2jde0691tOCyzo3n
AuVXgJ4CF6gRzEqT6NMuzqqo3qkzWcq5S5DNTxN4tsyzaclFcSijfribNuiY0AFF14MF1YIanOzU
q+kId1eiU2lVJyhUmPgls9oCIE1a6cDY1bpvy3ftSjn3nshjCIB9R/O1sSWCnYvhuW1bwNORgjoD
V0CzPQJG1nzH8hCMv4coLo6+OyNp0l63O1DgENcnDywhOxGhkI62YuG+hf2d4lLXf+ZcbXrk8j3I
6se+IZFbd57z2cfJZV9vB9CfVhEbWZ0xW8FtWlKL8Inn40U7UtVsFGgAuk7J1FFxaspstkK21kns
frQhGNQLiLzbS/lY9nrrsuokHCp7lri8c4QPCzMIfT08OlFHfYYOpBBs+Uk8iMCUjVk1DH/Ki9pq
erK6rcLZdGF8Oq3Zbkq257EmvCwk/l7KzqXxKup4L5pW2JI4d+GI0h46b+bB3AWfD28zKgu4jdl1
MhTaL+VDQypoVnUGaxs0+dfeMR8gOVwZeeQVY9ImfrVVmgRGJbyiuWWxFdP2tYJ1o5Kt16uw4j7Z
AjNne9+FXhLeGicTMxIObdHXDksZaZrJ3hMWb3kMVZczxH2QNQDdgv+avs54teOOZO6cLTABcTYr
HnIv9HtNdqeXB29Z9CaGKHkN2OoVNDmAOX/Eork5gtz8zLDuPzF99M/LwLPdmK4+TOTZjtA7VgsR
u5O3Nzk8fLgCMUt7+MgFlpd3VZDw4a0jGDSZ07W04psDZK/T+Umd6MpvnwU4vKhbpFO0MUfXgMgs
NdDfSy2cMjrjMfSnDbxUfTOdRpWSzajLuerjhht3kHFJfBVXsvBD0RBMYvPdo09ZsyUDtcTSDTFx
WyhfGU5pR1P8CRAVf4Uex15i471xOMKgjEV0rDRcd4ByBtS0rUuecNwHCIvJhm925TB5yBna9DIs
QOwPazSYs3h8NreRyQmsnTKT9iB5JF7OK8zT6E18CMntMr0hgeL2XlFlsq2z1boq8snbAHDCYmCI
4HJXmhxl03YW89e127DmmpvqnIMcEMwRs6jAplTTxK/E4mhPnMdscn1qpTsdfx19+0pcyGzj8WDO
eI69CBK7fpP2+jUpidLICi3hQshjrycxU7YfBCzKWyNLGYCHQirS6EKf4eVQwrh9fH5YO+t9ksch
ae4Epfq0VmmoYGUMsgOzTnpXyb+vJCOxFE7QKvRIm6GE04KRQB8xPq2sogBrFdpGL4mAJaLov1LT
rqCHzGPxW0EFwI/hcdADDKZwEUxQ4/rDN/akRpRVDj1SIQsAOIQHS3rm+UJAEFynfD/oPUGzpWZc
QJuscpLC4ICFVUnLJ7Qqe4hpEhkBYrUZXbKItSb/puH464Wh7wA0w17zlaM+A8RsPDW0eCvK7l+l
OXMse6B8+pFqY8gsqtE/icx5cEfJryP4voFSR3Gia3f8fpvp+y/Hx5uxoiPedCkCFhaZhzzUkV6J
JrGkuG564/VUisyCBWKbnDHUZLSpzrov9/43TrfJcpX42rXsMNHTdWJMod19XESvd0+oskS0yEJU
s9ml3znOIUjMehfpoE2KYsPzLcKeOKbHWqHgtf2yrsxMxOC8KqRZS8IofgWscXMw7C09e5XbhIIG
2m2Jnxcp/6ROWD65cb5Qi551qI3+WoePQtaXjVvn/3HARH6wupHgRGg23e8S48zsRfEbQ/lTZX9W
dp6gDWtLbXyoi8LVd/3GRnvc71ug7wLu2qHmjgKgcRg3ZRpt/iBUUbTHsBjYzkhYfS4ehGyT9hqS
7YXoJdjUG5hQ897l91hyANMCDcPIzGGpyO2Mk/czizNqgWo1hnhO5HP/fijvN4STytIajerBnQW5
/z+Qe/Z7jcZh82fbkJBo2B8JL90OfYfFcI+k6/by+2AeEj9gJhFOfWv1TcaXTKpQEsbnJO5HKKZw
cXbZ/zlX0mi8ZKeHNGFVbQNilXrUDTQ4h7kIILFi3LO5d/rJdagbyf0OJ0Tikqrch2lH7OyhfNta
COPAMom4jWB4AUPc8jY+4OVwjEnVyKyo3uaxcLhtqHt6Y579aqL+3zb+vfOTQwywmJp+RtDnibSf
tYDsCt36mIOTzbJfG5Ij8nbaPbqytSQtkzFKVx81tLqQKaFH6tAj/JAzkuaFNp80Q0YknGNu4+X/
tSfrWyMrGMFYJtB7jECuKriQw6P/yi3pzLkOwbJiYMGsH+MqLvL6AdDo5REJa68P9KpLRToQSFfV
jxcFpHfeZaLN7H+gC3EAaHYstxOe7I2lSaT+1KXatGPoUUXYX7/ZFoZt0oLQaI2K48BR0a6zzPek
D2zFrUfdTIGrohjKW0R1AUJCEcxst5dbQNwfzghEswAVhvRHgRwC+fFrtOqVXfd3DpWazLBnXAyF
NxZ84FQsiSRY+T2pkiGs5ONjlbR37nGSU6jXuHaSsB+6FUk4iUfhzGULwB99KPG9KQItmeWXYFqf
0IUUrja92/PNqyPSr/J+QulRZHwllD3A3KjOxsR4L7SnSuc7/7N2gAJ7rhp0nmm1vESsvEY18RNr
imorBxKkbQE6U/krWxxcKEKFqx8Iq6XOFKjJZssKP6EirE1SerETKoP5lpu72rntW3f3axUDIpf9
+cI2qmxACIG0Qjqg/CCluZzztAQA/Nm+yblj8gDi8gv2bHAk1MR8YZ3BwmQRA1R7PEPCIaOAi19q
1dq0ZskG7kptht3+oXQcZBaeIvRf6W/J5zyXfOuP7gc/t1DUbHmHx4C8DSxkBWZAfSOZEEwg5Qz0
pXPIx/UeFe4OXhIp1jCky5UHWqhi9FKrh1Szxr8NXMbD3rEJmvY3fD7gVoAgfT/L+LRFr7envEzK
psshvIwygeB7qLApeGFBaGRCYrgfCo44R7szDXswEBP4B/qhUJOq9P+NeS3M9hPv+SNqa7DV7A3M
LPwM7kuRAWHT/NSvjBsP8IB4/0bNeMG8RfR5vALzj+p2AObjKIptOVVNMblVXq4yruvtqud3e+KV
PIgD7MPGj8GY/7we5Urnljf4XWe4PCY0x/pVM3cjAu/afufNu/hbIjpQeciXiwnJgI5flVTIU3TY
Sm+d6ApYqy+3DJceHKAmF5zD0W1X7hy9W48Yn848L8AIG5LFgEV7ZPBgmrs3EVWjFtyuKE4dzatb
ifn+UEBoEoh/RlmM1KVwHXfDW7aqs8GhbgkDc/RgoKc5S+iFigOJfjbj7E8UpZGaysO6wgCgRmE2
FUTLPn20IbHhnFNlRr/cBLGsqEpC6MOcRnmp7470zIyyljzFJPIzDAQWmsh0EQ6dRqxA2P5zgXgO
n4uQhmtt19GGVVJbBdOQQEv1p+bsz4w0rS7CClfxLjF4fXUETuqXJMTwr/CCY85NLUDUji+FchpL
LWYthRULWdEKI/snWwdt8LTuOrH6Zq2WzYa0G5GmqBW89IB6hr6KHdCA8FrV972M5/6r5CNi4gSP
AwYyWOup3kDnIQ0LIFm5SoyzsfWpMwgTIj8gMjZ0xJwYoO9XgYzRpsOQP1kerkhySnVJ16234OMi
6UvXXDs7ZWKL7xX2N8d31eJynAURPbub/0S5Q1Tet0CQedf43yNpycjLci/I+GwEzRtrqMNG6O2s
sqmoBZZ7y/M1ekmiFEVYy0+Xc5Bcmgoh4qW4BoiD98XZABfYLHUm8xojBeuE0SQJwNtDVbS2dMaC
3pYOAYDcbC2GjEH+LpByrCPyNSYT2zOVDiA92VO9a1zKcPXyFL6uLxYWoPif2IaDm6LmzSsNExq7
6zRjNZe5WT9ZDVgizgpseFigojQbA+E93t9nR+wg9I/mkiW+uMmNwuYIKgfZuz8FWy8uOy67n2yP
TU3iQslotRE60PadtjoPPlo7lV3ud3MPXcrxANbN2b2q8/xS9awbs+Ja81Sf7W4yYyhaxSwRxipA
l3CKnZmh1rDwk1eCvG0cTb91EGyFXDFziu9w/bAs+9xECyiq+YevRzHlF6NLDduOTJUHXBS0iLOW
mDVJiChmJq119kxvf9WIMdIE7lFCNvOaSYwTjDgxR9k7iHfJ2PXP35gITcCCmKz/WLUFxiasGyvx
FartQFblRAGbDcThmItIAstQwLehIZps3GoTvcSUOYkKS0TGCS4JC5yhN00DtN+9LKv+YsVF+Nw+
6CAEzZNfHCv71xKtAZ5W0I8DWknqCk621KOURrXlN2sPtVNknoC/iuaDeyBEoIJ3ICr0phksGc86
7kMfmJ8uvDc6qQXdLnVf26hZkLV4e8bY8S1gAHi+lWPabzasS3Ah222l/cexpHaDgUenP08z+mC9
C/r98S+8D24NTws3+5mNPi4JsRzIGQ+SWomsRPKTC5VYfTgytmiK4PGCLWCemZuLG9EuhpOFQ7w8
glTYynpW7rSOYejQQPRmEkG1Omo7FiBthxWeIdL7svdk+gxlDjkr7FOCnqLU6SNhPDp72e3a1Hn7
wGk4Ry9gNE71UieNVznurqy3ZqlYQbdiTKCXUq66ir99NJRxMA6wHCoQtrEaPg5Vgmy4v68E9X8B
XnFJHrPjIQnkxkmVebewV6qOnDUH5qt/XhbdBMqB2YOsvtr7o2lLf5CG5u7DHAkDdZNJbEC+MYss
YJWwDSWkI7/UdbGY8KEQEO8aRWDl44ATlF2GfAmzEQYk1uYsi7LM58V1v7k6Isgwb2c3/8ydMnQm
3gjiDHR406Vxew6yZFnM5TBuduhIkqGDn+q+Ikd5XTigPpRJEc9Y2f6xoee3OVM/+YDrv0b42PLw
6jmy+chuPAHRXa7b6iFMliklhDSBBLnNOiAnWl71zPQE03f8S400JWMcuw7kMSwv0oUO7nDLTkhh
p8tunwUPEu+07UqIXRPAtyf5oI4YohLtctn/t34OKLVATHnss1HsIC9tY+lsAd98GFCJysFEAYa0
yYpkluPyPYUW6soxSpnXbeSPGh6FQU4sBtpOZl6hEmLQMfF1IVkCuig0jpHv6cXg5ttySC+fJ7UO
3clYhr0ZMaGUdmUN1KGNfJDC8PqJLZgNRd5yKoVrsdA6dQvp8uSUcq+RP2U9i99O9X5T98jzeA4W
Yjyk2gr5qzQgzVH2vrRDrfdUBmIVFHYpPAWZiXIFtoqsTZczJB6J3Yfa8eOsijd+VBBuZ8VjuuVh
N+9Dlfmq7pv9DVh0Ai6Wv5PvB3wwaJkrS7/40B5OAfmnxRtHxLyVtxgBTASMjXfg3EmqZKvy5AUg
n0IP0X+/cBEXME0NINnMCBd9c9tnj2xPqOKdQ9wErteghnm40rlHmg1bTw+TF3Lvy1cgyyxPVanz
CG8JB9shlhwWxqyD13GfQHNTSAPxoluchFUybGAkqT3JBTpOK0IWVxnN5aVyc62ch/bmj826zrTs
zyQ5710aqd1ExQYk+V9eSAsmcRXBS07wFwUJRMFW9LkK2SqG7WSTfzd4u5B0QIDrpvXl2VGhAbdJ
UEUii1OYvZlY0WX7vsKPCWR+t3wUaN13K2oORV9cZKbgorpvP28l3ARHe0TGfxdAUZVDu5Vu2APa
L0RPO0BMlFHC4V4UULly4gx8L5vNvyZYHN8Jtt+Bhj5GzznQIK8i3uHMccMSh2W7IWnES86S8Alf
671/kWFKRLFXqMrgt8fA7qCosO+BrDQeFz/UkMGbozHRBYvAwy5jC2t+RkLBCRwjsABNU3oWUCi/
nXL7LCbHVqGYwJJ1qMHJs21esddlrycnzFmnzfX1d81UWdjlvlq6oVi4Q3QV5ZndxPlKJ+EHPm6S
IbuRoM0+DncAL0OzgJdxRf4mFw+S/M+V4n/CCfPelGcwoCboSi0XmqlUh+xjcKmAQcmPPWdtORVD
n33v+e3YN3Cn/EhTb5pQegqAoG92QncKPKzBHOcyU8m6FCFfnB1SATq0E16+U9YNTIq6VMT3urpX
F6EDQDOQwMD237fNpZy/aYmqHAcyVXoCe6xvrcALQb3RUZtwpKWHGkC4MEvWnZx08vQjbqWnRf+w
GG5IDinaA3XcJ9DHHWatzhtRDcETpZdusK/Mlm3s44RIUu2WzylkNuUscrg8RXHctIrfeNz3hSJc
vRsuQTcXgjD3cyrD3KFnMvHsd2GDmXRVA4a92Cmn4Z9DvEW3XLgpf4rNGprU+ZZNjoPP1sj0oGsd
R7GB4vsNgQ1gfnXOHGY/Qp3XtibPZTpkqQ4Xv07Q8zy7C3wspR5lc96b1wA+Zz/uQzmk5GFN0aew
hQkJMY5rNNvXhoD3rsOKvgJVd2rardztIUsCfE1C5FWxUzecZuoKc+r55cpcWgDZd4AZJjFGMzdu
XZe3Wi35FY4n2osduVmsBk8VdUetoFnYOhAyUh8e+ZvIEdYVO5oHGD1jHqJ6ptapbPOlJYwCcM9S
hAvO/XkH8/hn4/KWJg30eP6vp0XbRjTnFdPM7+xXLJnmfeLZUWD4KfTDt6cvFdoqYOtgGNlcg+GU
fYdEKYC73kukHA0P7XNFjbECVV04HcsS8CgMM7ARSKaEZlj79Ybh5Mj0cmjeE0DP9UanCZa3yqNs
WO6IM+gjnspkMlsFp22ORyjpUV9ay21S1seaiQhD7BIak9cQ+V54ynzfpxKyHUbx5WFeQQYgg3oW
Pkfx659hLQWE+sBf+x7WM/OIXMV2sN6oIJo/aKIYVZjmGGlsWLOG42dERFd486U7wKj3DLB8LQ0A
2RcyixmX0h/ZycXAeiHd6eFhcdTgmMortwR7LQaC+nG4dy47TxGrLhdX64ofwlgKys6gbgujK1g5
eOaH3ATF6XnUftmL40wvdfTe3YSm1D/h6hvyuuhU8yl5xdXsU3pC2kTm9lj16MgYNLGJzvwBzQ7l
HQybmBaXG9k1vpXZY+jK65jO3k4nZsFG9hqjeH5fWTDaFE+n3EficKNK1VvDkVnf4KuMMNF4CEb4
8yw5SSu5E+bxWmcmrivfOR//L2bFcbPuCLBXGALjmCnmsBC4zzMNw7hecGTBbnoTBHGonsC3YOlu
tHybFduwy1/U66+wFkcNSNTTnaQAt9saWYocyIYDff2di7BnDCzFnfIslq16z5wAmdl6rpe0uyu6
v7pmFMu+BEsjN+5JEGr9+VKFjGTRZRiUUKYKbJVBewm04/yKU+i2tsGlNTR9wS1HXCkO0UG3q6RC
pZw52qZe1EyWJRyPCemzdz5kjoy0zW0jrzNFmQhwmZsa35+NAsFBa757Gqv8U+XkpzNS92+G2xtK
KKPhS1whsxP+NInr+5/RO1Mer8ybV5WZF/5Kjzco0DP2OOC4vghEw4+1vWYBqJC7q8Udt49oyOUf
3u9tFiyb6PMEZW1hgPMAByrBLd204DeqVUw4xgP8vty2dFfbuEQ4z7eww+swwTw5pyuwnH6KdlnO
LNg7Gi8jr4f12rmDyznDyLpsG2olVj6gr+KdeV6PgZ8530X62KV6XlnV6I9O+XtcS2qWXM96gzOg
G9Pa9MdBzZ459ZBF+3rYXH5oqg6gtSSpIaPWHA501ee5+SIwksUBVr8Uj3Kq+a4rkbzpml8KKJH5
2UFrrKoQ7jd0LbKUM05kY1j1f52SI3JLnfm8KdtLyu/OjLDmd+0lxBWEN7eEtByewzmYmIPa2Smz
lkdEr6uQlphj8ZfCZglmSr7oH8nRgsmrIFQU7w3iePUqiMDsxg16TNVUdEZbZopBwDWxvZNg5Naj
5DPCX2GDamqfLor5as5NxeRnrN/DrEaohNlKIp0/vV5jocSh8u5rA0qzWlouyfaVk3yIiWRiychE
XpMH5D988pEcChZIXDcqTi8cseViQBTROIMj4q4o5XFEcw3dSKzR+dRT76bYFpH36h1L79pHI0TX
gl5so6w0Hr/KN6IpwSeGfwaAEIEWDyKFl3/1Tm+RVJi85xcCBfi585uwYO9dhkI9vx8Tkcc2qggg
dfvTOxneWwFR6kCrPGuPze8wuxlX3U+sri/ZuTCZ9QPGgyShMw9vv+LgV74BCY9jWUcSKY+CZiTZ
A4h2+bJq7j7x5I9gEUIWdif6mJ8ASCoKIfvndsvsdWf7+J48mUHkCJTnRGEUlJxXCyT0ev/BEpL0
RpavdlCI/kadj7JF+bM/XhumL9+1UQoiFvV5FsdQiGnJo3aejysMtHhpU6x0FmIb7/tPQ/BcbiTM
tiZZ+OdxTiNekmRONoQVEPxJmXrONVkA3oJqnnHmt2ozcHCXNhHmZpqHfnf7f0TXG1hFQgP0QpRq
/HaWShBKMVCFi+czJQn/clHm5/cYL7tBno+tXhtLljS3+lM1ZJqDh39lNQglwYNirg/P7bQMqw8q
0TDxPgTHg1yu6FgsdKwXDow6cAdE6s/XolOs89Ok1rqeMmHnMvgfvvDYglq5BKFKQr+pYez7rEjn
JSv0BEc/DCWX/qYgbSQnO6iO7mP/K9zIAcOXtYngc6/wNgmQQW8gZSd0jRQSL3BxEVLlUMpxQN8V
npFzkBq/yWk1Jh7IT4StpomNAva/f0l1bQfDQktoScLJboqvKYDiRZ6z70VxdMDxQ3R6CI9D/8iI
ZBcwk+3zJ05gtLj/h06nWDocg0KJlOv97xVCdASFmGNB01ZrNObJCPDeBL1+NRo/u8C4w/Q38ADE
2OM4bD4UA1TS+rWK1JfYFInXKwyIMKLeFsMDhlQOWlNyfjNnPo8ZDI3lycFEn3QoTX8t9mC2y+PH
LJwkNl5Rlx+Ms5qc3YBiFUUG66qd++5aL9quT186vyfZX9u24Ll7e94TWrUKpEPFPuTj3c8Tmz1p
AGhm1+nhcdF4OwXGobjhCmNvN7PwQVoZWYGiSpd03wmF3i9DVwaPYY6Qrl8LaUAqGCg15r4cidwA
x/EoU9qCgq1T2LftPDwJ5WLYWSgcwd98pK5SJlJre4wW7aM04e7ek//nXhlnIiOMYS+EdlAM7OiP
b8qqRuI/qWRebwi1rnQms0pnYHmd8KfHptNO89BHVeuRwdsJj0/FFmfJZ2NYInpE0M3suNpNJnM7
j5h2PDs/vWdPRI2D6V8mz54DLo22zxKAjgTeVyYWDxE8s0ROX8QJDqXr3LU8HVCRQNVqsjZwaIsI
d+ZSHEGfiNGIC1brsraAsHscVVqfC7ksv4NK3UkkxwpL/SQfPUxTDZ4J7mNES8aC8uJf9/BQeMr9
dzqUIon1n8h/ltYWtNWqOZIvWw7K4Uuww1FXF4OBS20+Zedjt1Q1hhANxZTNwEGFybTtMHcipBhD
TPm7HWt0DwqQdKMLom2TJyiM7diQMeUiWVWHYvl9pO17sS2EGq2pLBhnNtGPNuZ+ZCAdESMRIuPy
NMVoPxxdXWjJVZqBR+ffJMwWl/lRhJwU3p8okNv1l3Okvk4bpgedxVL+Sn9btjIRnG88sjT9xaRL
fAwUFO4wu/E8TE7nlLtjtLFbGHR2uVxlKyfmRxvNUiRI/JOYntiv9izhlZP1CPey2nN6udIu6jBI
vBufkLD472ceQMhipPAYGn6x1H489N8lU13EQ+fbYilSHR1eAk+CL/rOfh2fMKueDDhPmoXrks4r
iDb5ePJ9f5Yyq3aZCMHNfw5vY6znRqm3/CLRj2qLcYZcpDbD3m6U3GXph9JoWvnbT+q6aeywoduL
bukocnf78j/ty7T0Acjeke6v8Z+Yaid62HZ3q+/hPBRSti8MG6My/rHraNbMM0DQBtWwKyPtITia
dOAQTyDO88Vp9oHE54KZ2RP+xvi3Q/YFuTzIG2rT+hXWATXte90VQRhcbayUIqA24vjcvJjf5mMr
K/FbjxAQZQkuVMCMAiGHntN33J1Ak/nlNmVTgMRsbnl124n47U6wRIHYta4e4XVhjSwQXpsPRPNE
AFQKuOMzjAVLPW/6E85cdzAac4jtaDpppirw45RY1fdbiEPUgdGxsuf88yKGhAZWqg+w1MlGgzUy
PxxkjupFHfTMkVfjTw2EBrZVxzLn8VzWX16ma10ZUyCO1vMuW1MSG8PZpPailrrdwq/f/Lpgr4S/
gyA6AEXBvhWdvXcWLhfYSQ1wvrTe9GkmCjLSwBEwZL2wqYS2jng8DGHklolEpY2Ss2+99qTTYrxZ
xku9+toxXC37uQA9p7YkgvlEcwhtfwYZI6rYZeKGt73Wx8aXZlszql3Xn5uZ9J/CkaHh/Y6Y8AlG
zxfBNPVKBuJph8dCY9Ke5uj3U8kl3FRJLewACEc/yJFsvtuAiVrxNGIAOhqkuEbzdgyJwHujED0H
XxGYLdgQX1qqoQAOQ64OAydugQsk1TdnuAgbLoKWZyRg8QBnY6YMCBNdregS1mzT3X/YyFjo6sJI
GCKVhos40MG9e/uTZM5Ab7FlqpRWcsIR30sRgMQaHMvA7fpU/mken9O9LyPMtWy6aD3pULTfEOPw
37uhhWjD5I8HW3H99JLZUAbbsBZQGIlr6V054AujdlR5DInJff9JVqeVTyIDXbeUzawwilJ/uBvy
eNeKmWh7sm9PVL0VhV3zefJfMIxpGaQLt4ohcnkE4CGReul+lAUs7VUrrh3PCea1s5B87cq6jhlT
6ChkM+iAM5qp4UnY04nsnSeryuW9+/6BROvK5fTxF+T0StpKIx7Un/BX0vJ6BigQ/pcUmQAEmBKG
fGpovK8LzcQPg7J2ZmiD8OYZXAt6wBaDTDor/zCS10NZPEAWK8T9HhtGvCpxur7sxTG751bWSZ5f
FqTNNkQimVUoSaD7eZQFoJLpRh15FZYmnCvPzh3vPtLbI8wfhnmd7H6r3670aRs6WiRJnQlfJC4i
RrV350F6xxhJSMhzilgNCzIPy1cQ9ZIaRyxYcNk05vq76ZKh/V3Dn1sRBBzy+R+F/5FbKozz5yoX
mVQfMMAsvjD7ic0ues7svWKI7O7/op6CWtGHu8ZyALWy4/HEQ1N/TyA3cup7mxOOtTGE+XeL4E29
Kt4JEdHCsuQxAfNi15aJ9wEWZc4JpvXLQ4CnRy/9rU5J48rGEQtxt8c6INSjhlo7EawciD6xOHDE
XDw0tHxRoYP0nJWtl+w6l+XkK1JvVJbbrVPoLmjeHQmH5O+PBubFqYsHrBiQ+5rPP5CN+MqfsGLf
G4uOSq6hRRWQRkh+ZP/DuwWVHuVCmOZeR9+hxMLOOkGVTyQb/YSjFWFY5nAUbKEIYjDvFqjSCMzP
Z98YA0dkQoO4Egn7VcYChjP40F9U63z1Vvy7UDGYTnHKVuB6RqmWG6Yzywh2Vwa/ecpjM4sBxwya
KG6KnodWDQPe9XjLupTQLMCyDMka597AeqF6XZO0EKnpPNLV5de//+t8hBE2QCQ2lGr6jYfmdPBQ
deWa7O7oXsPS2ekEqhTlxFX18LR9rlN8bABdJaGNvwUXABq04v9rSizFHHxkcIP4qemrDD2jChKs
m492omjktXvzwy4v4obz2qdUUjuWxNehg2vWGaZDj7CT6Vqs/5o5VWYFoXGL++OOUINuSUWFueWf
QprEkzandMGtXvvsvBAuFFpCGENuIoCvems3wFaROvkHWZk5Mp0SW0AYsnP3tN9PzcoXO0sIdIDF
Gcbt7rZD02WEcP0Y1P8FAJXWg6Vv62aqSBlq69fhFJzznhKtbijlKKaHVLlKu4mzzVWQiwIlzwxI
lLySdD5Trdwod7Fu9tdsvoFZuvu0lyl8BZ5oY3Ix58D4g6XsRX9DkzRrIHkxLS0S+ex1oboBSiiY
9haF0Gkj6kA2CXWufRVSjdc2pQdoiIxVgVXi68jGLe4bc1+Vvhuc1YeWf+3mQCOAwRpL8HzqH7/w
ZXdJgEsyceUc5uAflOw2z9xZhm2uBOBs43EVJo+sj+49sF4xsc7HjVAr2mGlkwkFk4327UkwcHwj
hsHS4uR1X7dzlzkyS5WX9UCqKFXHM8/LKp8ZGV4Yio/meQzeE+9gZRjRK63bC2qC5IDA4f0jwRh+
B4/gu6lkTU+B+T92nxFMD/ewWaKSH3cie0jP7IXuBD/M/FBQzvz9MDnGWTde1SX6c0/193EenSfD
CgNqukOsHjKL05zCVrZpXCs5Is4Dlg6d7cxgSQT42HvSBeiRjQCqx/Ws//J79nmgWSm1Ymt39f6N
cLW3sSZbADlZJqSCkL9GGQNkKe+az1IcHRgELmkW7BjGTqj+q1ZZbZiLLNklu7j7YBXYe3Gic7Tw
NEAz5Yw32Nm7UhNxjg593i4SdxH/mergKeajK5LcpXvqUN6WfGRMVJuXcFukNs38e9lh8Cl/ePJX
RKME+P8+FfjfuoEWayq2nEcOmv6HbFjFBzCSQ8HSU9YXvpZgiyWUg+bwgToyNIIZUufHyrVBP/0u
STx5hTWoVlGYeWOKrWA6D+wEYHOXB6I/X8bbjd7pCqNEXlla7zNyWn79lT/1qciJAWqnr2ywS1Bs
k+HPu/4sbsg+TiL187G0aYr7jOWzbR4CycRgo0SNck28x80Z7Kp5VV8vG1QbCgLBHneMWFw6Re1X
2jDGgVv2WuxSu1ajnSGfH7wZumSLxGyKudJBx1JVJ1sZI5F7yA1km3rJkv04gbU3JwG0x8rq7VGg
yNNEfWD4/9lSX5vnbVP3MG30PV3+KNAYaYEldx8z0Jb9/I7/5UOUmhc/uo4twHWfl7i39WClHVlT
bsmVqEcz/yMjV5tXUmORUFgQaUCU1xEMxtDqYuLL7skPt9Ia4T1tK546k2FZnXRangAaKxM0Ak7a
1HowJnhGQWUfWUxs7xWmWo5DVnFdLQ19Jkl+/pvh69I4OT8IBb9zp4U+IiuPKLBiSc24qO/K4j49
ie4sgaPS1xKJeWqIRzQnYjCX/3e4z7OeZmb4p2iiaV+5I6j1w0B4u//1WMR/sEzaGD7wT8Suj3ZI
aN/2umk1ydoAxPS0cLDSYQwinvvXnED4wovukwHc0uXAUShYA+K5LeWReNQa5IypsYzWmhfDvakQ
ovuX2HNFXrYRDZ6ytLUjOJPfQOVDG12/znTdSTh1geZ12Vt5Sep3Jqq2YhyJwEl3Cnd1K+YHx94C
GsMmNjOimkEkQbHDcgImgReryzUxAsABcbhW5bk75mf21E9KxrRqlCjrJG2/9+J1y/WOsoJLKn41
zKNeU7upLs84nhup9nPjmK0ZYqtV+v7VwmVxz3aL7IQXFEZS9qOHpHNvDMGme3oJCUW8qIeo5Wei
x/mQN2n1aK5ZeVVSfk6mbD3zNMqLB3MIUYyg7herLnhwx9Vt5G643gcDueabSbgLlJqLOHMmK49d
UV228X8IZMfimegzCFnFxNetCwaH86D6wBDPEbNciRCDfqfvpt4+P8nCZEKsBOVk8k0bbO2sZYmO
N9bOdT8UKZg35KIB61VwPTBJS8JYahHQXwhYtZucagxeMyp04aMB//62pyx7FEh6yweVzijf5ZO3
cvoXHoFARC+RJGEzAYodBiLjoavgNEjbnI32suQmzJ4zb0j/OF2imesUYz8S2NZRN/ZOZh/cNCOc
0SP1K0Rt9Xt080IJrR3LSsO8m0f7XJgmn5BxdMglfrG6tJ7+bJjPi7OIGUdkIZ7pLJfZrQjs7rEX
wVizE3tdtGfHndrMcWZLKifqLUL8a6+1YjD0ZlyWs3hosuvQHjzeYGB5KpnZX/D61ufPEawYpw2Y
2TPqGh0jHhkOZF8RE7AfJ4nS/khwUixLtGww5UQ/v5oZ1lWkn/kLwBzJMDcBwG+gPF6GaacejEOB
GayIMDsYMe0nRi6PhE9OZldHAt1czGtRjixUEfHhlRAsbW/Xb+LpoO/lxsapTxCPtLqeEwKFgf9+
wV52zx2lUaK8mHuRKlshoqhBZrBt9JdNwaLt/InOZCGr7/eQeAzS/hMfW7EK6zSLGJ+cod+Um3Py
zhDVHP7C5gj/08KVD/jJPLDSbIq3079YYH3NJjQw6TiY02YeZ9kvdeUu8pRnRhwClu6Zq6W38b4S
2AFShW4NlSYhquoBassX+axQc869qhkPumjuvja/mKEqLyc2/6WyJ43jjq9EXU1lQ60psc8WZf84
eYe9gWvUoaAfi4ENMqFQVKbZeKOPqIQAsR7F0qNCiLEFn2IXGe5nTGdjDPpqcVTUa4Vb8fcleSub
2SKzxvXcKh4M16BJhpiZebU0I6bPU1cgTuLWxjJrUwBatm9aiPhmxKETRhEBsUbByUqPaG7KCMSE
+DcOlgxRXzjRokEfpN1H8bePe8LI5yeHUYhJR7CqSShNkV2XVM84U1wZZRwOYYn2tH6VzS6DUgaa
gzgWtyz6tmsyf1q5b2OeifHefxN4RV5MUybnPjW7X9Oe+dkmwo3ylxcDrFfSL3q5mtZMcT1VlLPG
dczD+GrMCMjAE3urQun09W0XCL4JYIGh1dPVyWGQxhrdAOLUObZ0x8jY3ZOKqqnl+TrbqkIVSSBi
q0I0bzokdgldz0yPfn+nUAlAcVPxl2AqQP/QhE7F7pVLue+haBV/q2ImHPLSbe9NjJaphZbqPcrL
ZIQVGljHefmzSeuWOVGv08zrW9IjIRxVd+1sTxYnormKS1D/g0uORe9D/0yZoF+96Uids/lILsSD
kbhzuCNvXi7uJyjE84NmAitoNGbPQQ+YRQqdGe+ErZGylU7y8dl6k/IEpFWnA6ZlJvi+fVGQFZ8J
zsOtuzLLl9WgPqHsVSVrURRFXuneTcweXHKnMrjtiXRi46Y0UDQbyXOwreixXadgmZ+8ZCC2JXfX
37tes5ag32EwJjrc4UrmuYE0erHWbMHLZNZKdO5W8F+6TWsD6SHXXH6PScmcrvTNNr9y2CgbKazi
gXCjl6r/dpTIjFjsuwhXrUgmRzhc0zXchkIPoi1zcKh+0z4f013spbe7wjraLBqnR8XU5KLsr6/K
W7Usm7Kls5XmWUqWyV/ZI8suw5O45AoqsqWThhZCJn3M4Jbg1PEPwRYzSSTA2aGSDjSCA8YSpVxp
LwWXEB66kjq2wlfqJttarENECQXWbornNQD9zvuibN1xM9kDyhA8cBGnB+PKGuByYBSYWW1YxR13
reyIaIf6de9v7QlGsW4Q6eH9A2pJm8VdtCufWSxl8gRb+CTENC8ic8lgiIu1zlk4Fc1VVNvnLPg1
nhwHFk1XjsjG+059aUcWiUx6kjRVghVgdIFrdUcwDxBCM00C3WBSm8JBKzZADwkJeBtkdUrnj4xC
7N95bdNbuC1nz10HfPzKS6AlnUzLYlpsN0BHSmXoSqW/bCxQYjnvXEpDydAMQI31aUpxWcsvyyMQ
NYLVdl7z7FEDEixtTEmUvnKMlOEXiuhzhYXvDxBKJdI7m1JC8etotEP8g/kV3ElgtjTrNFgJ/KsR
2TA/XTaddGTVvMGE5bq+fkzV/ohY4qnt2bvXMbIUVoiB/ALtKkYwmlZvQ3bPcZ8UEolEed5Cn9ma
GVQ6LlLlKpugkRVXz0Yj1tgtTnf4C3w0EsvYQ04qiOPGY8iXiavVP2hS3jFvFOjZL3P/LOjQm0EP
m/5skF2aCRjUpNAvqfAS+7XQQ59iFHYkjOtyHeBRImuvif5ANl3DLsjgNMUIuKMivArj+YITGVER
q+dWHiHjYHUyorqIHiG2/FfSdquCL2rZ5th5d0Jvf4AQC0OGszMRkxHNQz/JXL5AFT5c3iBfqzvq
S4ktd6ebHXF3jzfqefPQvQhOpFtCaL/wZB6eP78U51XW3jkizB6pwjeKWBMlQRLtVcYF9+AqrKY9
J5TzGclBAd30BP+HSsI41Xf0O4NhsQ/evR594+JGiRDNgfT7OWF4GE1Qa+1CykQMKhpkpKDXx/u4
dzdNWbiQfE2gC3EfditYndm5hXk3OpmGOH46r+vPlAL8JNDhmYvkRh3J7wHlGbNNrG/qatoLbTCY
vaNkOdb/2Sy1r9JMMz8t5lN6YitHYT4DIkL9B6DLE/W2LtGu09ixdtVvRgw/2zLslCD6XVGoIGkW
iDxTyNtOQdIRA7+NW+vMeInHLI2J2VFPNaalF8YSi67n7QcV+WXi9iEm8T1XYoLJMlkAXF48Tx+a
b/snPH1j4rF5sdHha8sDSlW6p/+VyBwItksgbbUufAQdc1wxdz5GjjtDfbYgtb4fWakoSikzNn1D
KTJraVih4fmIbjUJ2F8fcP/fteQkg70AVgPq7OiWvYzjh04cGjFrlLitBgB5JgDPvTQphTK74+Fa
uLdcwru/Jxvo9ZUpeQQ/lVF7Ax5CMIPGCwIHYrHXWE8YxSAdTH5kGhw6/7HdbYtob1QLiYsuOC50
SXEtVQFMtl3lAh4LV/aU/1Bv6RHta+zhl/F2fmLmV/HGyvZlRCDllilEKmJc4hpvXCKy5Jlr1vHw
UDRjpotOownrBqRss89ZkREHzS8YHE3cwJlmb4oeUXxAzvJshE4TA6uchjScdkmNRojvAH2f+LBQ
OyxbvyWMUBrru5jB7hnTUnf/eh+BoLQ/TOlDENRE8/IcOepAsQ/13++uKiAo4CGOTS+dfPp/PTN1
Gselhu2kE2mBFBbBykvP5xXeaUXY+A7/nLOXL1Xyx30XZFSbE0zrQL6WA2xy9uwA/UXn7VPpZz8D
RMpf/J74hcN0Cxpa2sAJYza8iStp/vCrkvBwBKuA5+83pVsv7uyHx3yCzh8ghwxjMBdEMygvjE+W
bmaNE3CJyH3IOLRTL8leJ8eUYdw5go/UsHryupMMuV9o/ROtfaj5eoMuHGeix/SxhviOCTZ9LRI4
+vFyo/ExbhKnnToJloGBgLJzZJ0Pq+lXUKO3USZwPsy56gKpSj2KqPIpP1ccVnxeW1TU4PmMUJq4
+46jjQ+XTAbqdwOPIEd4E6S6+e0QOsEcsLSxwyqSEmS6WBY0rpDYdJFPTcWH97JsHBR8DNwwrOXr
8avlnhrfxPVxBmQsZNHb2OMxAHEsuu1mifsYohmBs3CId5bkTy4GHQejawv2Ay8Ms2C1grpkqWW0
/D0vDchcJhz/EPH6Q5f1X9Hf+6qJa1buvoXdn9RbW3P0ipMJDLzxTWfO3UxYdSMcr0//zEWthyWu
MIiMCK9U+/UBgtncrCXI/IxjFZfTrlt/NZsTPkgEPI/OTxqaOE5CmB5UPywdEniQHd8gRPM4GGOi
WIDQnPQSmXWaPnQWFAk+Ol9dIaT7e/2ufmYReoDP8kv8WT7PYqnueyo6abChz1ElI5qCkflN+AjH
GY6dn3AzzyyG3csiBAn+CiIjyWUkQFBSKdSUCq7T92G7zZcjMoqA02A+lTov4LLEWKXh7pIsFUjy
eVB08ViT6YUFJBf/0VBMAxQNB5Z1K6ehNQBw/3XICPTREmS3eFBUVMx0mYQNOG4jWild4PleUWJR
9OtrCWfxzi8RkB7ERb69YZUMi07pQGcn0QLAxOL+sOFpLkd4nThIFr3tdUJjukLLMW9vW0o9jPrg
7IAaIDeh6Zfa8eV2wrTUu3LYQDyBJsxKIuyorAe4CuTRvv4yiXtmEdWUrO1d60bCE1nCovK1wNoo
SdRistWuduX4NJtrwYNszhdWGm7Nt+thzN8XdF75T5JOlBSYUNe1exFuS3QilyATZwwz9kxe5QbO
2ETgCktSRIUhpC1WUlBF4pxK0k8MF6/QbYnfswCl+y+g7Cwcg9n1lVOIy6u/gAA3rxrSEnp5/K1Q
ze0Vpwpuq9oU/rYyuFspxljS7Q8zKZiifYU7V4B47F5D7B2S/qSG0VwYIlAy006MAvEy/nvCLICR
Joiei7eltaH58jG1UWEAVAFF6VqSqcA/DddTUqyGR1fIboe6IDqfcsdZPRHu62MrXR6mn9/n31OF
MGjMNy4NydXpJ2rEfGsHV3Bw9anVcFJ+LhAX6gi3mEUvwFm26MX3TSanfX9ZO3ycw35oLXBQqh1F
M4QsGQZ39hhlJ/TKcxrLKm/QLIgXvmOl+1LAVrTK93Yb/4+1xXnHhxp/2jX/NQCr0/9NmKOWWph2
Z+WORhWerTV/r760ITupL+LSTcVIGbdDP//Q6HQAp0PREuu3USY6rBV0iROXdsRgK5FwTgzcxOyj
IGuf/t2R0wcoQbChQTKFn9LcDTj2q/y9fu5PVvtSVisWbJ18amqsWH/Hjb6Z1Lymje5eU8cQybvF
6JLHvLi8/NGxSe7EV+6gIstfqf93JIFhRUwP1lGCBHPBsQTX7c1t8CLTp2yvjz1jK6fJOSwdO0Q3
XmrVaW9hPTsjOLIst6qRXgVw2URFT6BwB25wacoT1MA0oxJBzqBqA2WFdxqk2J6/5v4ZvTUmyyY4
9SMnoF+ainggwdCCa4Z0j4DtaYj00KsT4MmmXMtN+5CleB7cdHviVF+mruClbKa+eFtYJ7x+EtM5
YHMcBjigjzrvk5uFqycUmRKVk5mXdeTrL9/ZqKdb1jgYfE0B5beNLoEF6d0ucfw1+EIOMvzaliVp
Hh3qg/kTwDqp7P7Mzw0XpJLY2ZwWcMBSZ+lUURX8AQLrCMmQJ9yBXq1BxmlQGDaTOUJLw/glRrrf
9uU55d6hc4Ho4l+7n3OUWmG+6koACuZ+CTXb2owhkzNRYeuXswdBI+P7rlKU9KqI0j/8tajlYuJw
Sy7Y2iBvXWOPkKty0B3GUs/9q0ZSg/6bNVSCHpVIwS+Oz/Op8oUfWWR1TgzoS6y5/lQcfhHQgTkn
SNgzlmku9RiBI7XdnJJqtZKHx1TkoBHfHKsrUTnwnz5PWzks4etLFDpJwobucI4K3/u/sjBYPKSp
56Evpl3lcxmOpXx+IMTWuMEWtXm4U5iaDmhvUhsDnrIgytBWlynRYbFTsn69oEpmY68KopVSl29q
2+geGGzHfSb+09d00g0qquCxe9AkMCSwKN9KXgsaLPIV0DS3NbpFZEq7nbBmEuSEflsjSnX9O/sZ
XuZvCdYYKkgTeaOJl3JQM56/ziI0aKbNf/1DIcE2/72s3yM+dmwK+aS74TdlJlC0R4oA0et1w3xS
+BedlpuMVjmoFLfKk86FzMx8nDAszh11visUbKqiTj+tA5kS010c8GUYY6Enc9WLzHWuUjKDQuKQ
HGEoZin312JThFg5C/CqitBTbr0NmUjDLCphSJriOeq5wrKQI4eNyGbqEkKpcA9QdHMr/Jxp07Hk
K9iJgopDnRU+UUa5Rd92wIvcVxuc7rzJAR3GO0yQLxfhK6dgEApPzlBkvGy9a9gKq8X4S5loF19j
u9Fb/i/E1qBjGBLOoH6ykVA2Kg8TOiElcDkPV/Wk93xFJbHsg9ZMXwteMUIYv0JgwDtponhze3l1
BRHK/w6Ck7iZznXPoHCbRMUgn6AuksYt7BzoRsc/hMnjbdnvUgNsf4Asg++51JtHp4hjL4c5HVZM
VkcH7XNnVQ5rx4a/tAcuLgvxk3H+Ljlximh3FKwT8+8e3bjZ02C0SHhILXfVIFK1/sY23oGSB0ZJ
y60uyAN/8XjC8qnuPnCNgjhRByhfZEGyFyJDaUdA7yDMwtzzaZ67jRgdiY5GYhXbthjum5bQDaLG
DM0TQ9tffWAAkgQiP4YjnicaLsWaJXimvGzxY7sFDwe3sNKg6lFnFCegYasOVlsIL/UUiQkfOIiG
JhcC+Gow1ahoulqc+cw3P+yNjQiIJLdGTH/fK8CdRhRQlYU5VtVKzjKUfldwqPWbU39PMb+7uThI
lNn9SZlzfKs8DFGUiP+2v/jNWAk09C3pJAbKrkABofAqDAJ/jjdr2onjDNm/Tr4F5jTQQYJCZ13R
nThoyrjB4z1pAPk0o1Vus0qtA9p5orwPBZuqhnXD38IUS6EaIiShY7gmlFQLvVzkHUqsmMRVpxbi
9PicXry4LPBEJ9NrNDcUV/TmY9GHD7uGKuz0tZgRUJ19vrYkdaZAbuH4Bm3wAMCNkHOCaHHrZYLH
XqV/QZVE5v765Y1yRFjaDzNp+5s4GY25YMSfvp1h+wN5+rt4MsfRsXefX+ArbdNe7V8CKd42We8s
n1cEPi1lM9Qbcjt4zJ6Q2cIEkpgA1eljVb9WdKI6/t5F3xKKj1abg2XOYuxG4QTtAejbmwUjdknc
YNQz1Pvs3dihJ6jQ1klkwwkao98Jfmx7i/T4U+YNgZygqU4KKocVapxxXaSVVScPyxAoq7HryIG/
ip3qyIunEDaLVCogep3cnPjz/fY+3mN4Wx4Apjr1kgdZ2VO3InyTwKrj39byPBFOOF8e+2SZWhWV
y0UAQUBKCqwdt3xpyxP6xo4qgbtPSDbI36zXvGu5T1B1lfqRhkKfb+q3NFohjW+cLxryjLIQL//M
eYY5DSqqVBzcv0Qxn0FUCTFn8kEfpEp36p/z4nATO2eGBzLzR5sQ949LoC6cOCSAlPldCiCBV0N8
Au0/a+34hrQtMxi/YLHhno6lYZoeYN2moUIRMqBSV8UCwuEEy2XISoLqLhV6hdYtX8AowVsTYv1x
cTSDoIApMlnONYlJSIEkpvmd4sM6qYkeOkvCEztf1cIoa5DW4RtOnq8058qChdrqoVv+xiKYQHNH
Tg5wEDttReqhsDgKZx1/LGU8UHtQVHluWmQVENzfHrwuEwd9yQlcCXSlZNc9RU+A6CHuImDTTVxR
VZEKwrLlycGponTRatyo2OYZtLBW6tr38tayzouPB7hv9ng0s+tUtGqM0fnjfEr+gdLzyP0kVhNG
5jy13BoQZAWASjwL33jaHo1+4Y+PurvfrqCMKiKM3KKHS+YzbPP6B4l8FH7L2Qg9bfZmSEac6999
zXTNg3n++90J5tjk3tqtpPp+8x+x0+L2Etp9bSa6RZkxi6RILTS8oLD919cda1JjcFcJehUIDA6Q
WayZdPeimXvpFJxtJFPaeC7kv3rHI9Y7okJTB0P36z1P3x9mtN7l75awn1SOLG6bF/ulVH4Pqzob
jzZBXRmm2FxEfOOWBqx+vkDukICD91yLMOmM+e4W13/iP9WtzGw1DuDxKxT7BMYqMsYNScbxoM3s
8BfUPwhS5Zb4vlxwxUwNtyeL3AECI7+qG/+vVKFYCdfn35n2IDs69ryuaWTo8IqpIJju9xTIDKaE
tJBcCwc+mJP2hwthD7jFahhuM5pn7gyffASw9x4l/dkjbSs2AdVvn+eZ6dRLP6sMKhEK1lHwAQgR
Mcc7Q82uM9QIDaIl7QLIcfIElYcOYDzUIgP4o9wLvkmUeCx7eetl6wu7Qn/MTlwlf1We7LM2puPo
G48wbE8PHzLRr0czBKrGPgYRk1EBloKIs6+aSTdUH1WVDs+eJeI92JBbFFfTrIIWUWIfAzNnHajp
HL7N4C5EXNo3ax1ELerKLHGSlWVQLlSY9vyApn8tUi0wdEEB1sipNbCX2y2h3QgXDznsWl6BWgex
oDe7u2Rk06KEolUgleK17qA8Fl0uBH+TTDyUXkzhk6HhVC4ar8j/NbiXnDHqyq+cll3YwJjDn89m
uS64k1e/Is7iRcNZsJxNvhp+Wdz7gP/4kVeV09ELx9QzP6EaUMclFxC5O9GPsYisY3u1Q0JD4o/y
0PpiHp3yHZ9RXbTN9hosRJ0SGwv9VvYCVLEh8FaXCuo8uML0DApyiKL5BhX78MAMhggZXiMIV0rB
s8+R2gTrqxP2vA7e0LsMJtmFMaFVIGjISCN1HgjCOmmhBqJbjc68tgF/Vpbqhenc70dUUu5R4YF9
ODfXc0uaiOZDBlI7xF/6cmNSbv66kDRlgkHhRovsH6KqC5IpSaXEz3jruAfizHjmGEl3wm37csVX
B7tfZ+iRsg+G+F2jxS7E8pjfn5rOPRZ6Sx4LLk+NW3bDWyxS1Z/nJS5X4bBwARk1BuFjkp9DpY3x
IMOahtRPwfGC2f9pJ6t8Sv2RdcYQKOrpf0kDPYXhqiHjXaZNLa9u1vT/UPtylyHz+3W7FOUf1VQ0
qMoWs5RQSLBtnxZSpOiN38p9GjmiKY+RPJHpa8hs5HsDJP5cu4IS6cdXHZtY6f/DpfPMV0v/ERNZ
llvCjgJKWC8ESEuf9/D8/Hid00HWAeB8293h/FE51FOYi93WUOS0ogIvuXrRI4AGTVAjF5frMq0A
faahSbpWx/aJC/1/2uTNRyIcaH5Cgs1KaSn9u8zu+ksECizL9nVOK3uUqOHWSDqeO3Jy+TIbtH4l
4bOvQqa9Ayc8ndMlvS6zAfv2awwBsWYznjwa0ekS65S4hPNTk+MUw2ib3D/hMsH32CCABHjk+/ES
Wz25I2QoRs12NlydZ+NknZG3LBVHp7+RG5ioOExqA4bK1eolU0QOCzjbppX9TI5CFYVJ4/HlHFRV
1yod3nPDeCOxNn5t0Bq4Uke1UhHo6tx7wMwkLSSdorF2NRNdbkHyF2yztEIbOmQ+Dc4XxZ7Qemox
V13dqh45vFK2jEV7b6iX+5FB8oNu8mfif2hAp16zi8e17XIZagPf7Faf9RoBBgt3btKTCatFWNs5
0Zubx84IywkTt0+q4TZCOGCb3G6oY54ed3sWD+QXNpHznMhpdD96PjcyGxdStX90Mdq8WhtOVM+3
v6viCj6+mRapyjEqTfquZMVcvHpjyJQw/AxVpNR0DBMgf1puO/R7RZyTe2cAp1tPqV8thDb7MOFm
JBuSoapd7lAluW2F0eAtTy3Wkd2/fdjLH73iY8UO8JlBwE+QML0VVS1YaGccLnDUVK03YNIhE/iE
8dKD9G7G2IwdjRvDt8u80SlrRUCBFPBbwL1ke3la9i3hL5CZUz6V8YUXno11UeKAZgr5kHzRyjt4
u7smTuw/GHdZ4KYUQBicaRqfQJSrCjynHUn9i7eC9gcjLbFoY3n8H9Q3Flo3KdB6diLFL+KMczce
Huq64yoD5vqNDxfkWNauFBGrS44soXY9CP3CjAqfQoCs0xZtGi/D0A7h/tCbfuwe4aHt2U0ar4W6
fz5FhHc6yCQrPcYa+On4+9svZ3W4xu/EFo/l+YCkAUrxvGZK24FQf12nC7W4gc0/9sEsDiqfSiNI
k45v6mpKs0fFPwzYs9kfvljeMaOJBC6uP0NKlpsRh5pBR+xXfUcnpLJinwLZ4u+bOir/fO81k90+
DSlcjIYzBZRvQcKbeh827f58sBXDr9WYCFi+Sb8rFx0kp+Sf+taA+BaueRYr0FhRBeZzRYOAHG/W
OasFdhZg55JGeH7k0bD0k6SFY8S7Rk6sjbg6SkPwqb1+sEIDI76zHdsEnKTLX+s7Kk2GseSyzW/p
k+PiFiqLtzjqk+xT5sgwCQkt2NoA5bjMqpw1nvFX+6ait4rqz/+TpEpn+AkePpAKiOfuFVudzo3C
sBpQAHPpFsxc1SSPDE8OJ1LOTqQvPaKojucCnDjKbcCUSx1Civ+Je4B+qFvdjcZHumb9nGX+qiVy
xu3qXSOzccQRHALYG+KO9LiJqPr4i9gl8mV4GT07LJlTHBCjSopgUnwtoldm7MI5pDXHnOvBstXb
OEDyG9jPqnLT/xhGtAQ4q8RV2oRQMUN7BiqMP01BbxKNdzuVprVS5FtVTSwRaB1JFMPMyLPMgt44
U3zc3hwuBJYDx4bQZHBsULUwcFozwofF9DEm8tRNOU7aQtL2GLG4KEoCpAFwZEnJgIgdoBKWc+NP
1ijL9a+GCjaYPXasAV/ttwTwPWwPhlFrV0bEIQUGp8zReJYenqZU65vprrcElarqQL72+yaEpVjE
kIocbAcZ1A9ClDJmk912sYtnbopSjOu84I25tKQ2wUgJKezuCXt7SI1DePB8svKAmLAuG6XA0Qg1
foa1dIF8nHPdRO3mRMcVithos5qTapxWu4AcjLmULMWH8WS0ODMkRmh+/m+tG0Kub9rvbHXRMR1C
wGQJBBLeSt1vHGHsZ7d3SSsR4A5cpsDW9kMmfTRzJFUz4nfTB9VMWTcaoDL1V2xyZ0AFhdMiGkV6
HgoTOsq1edtou7s3YhWZfNYZieSImLOsgTIZ3+XRqNsn/9a1ZHdf44il+klxaoPhbX17FsusSqhk
V0S84ZPWoP+aPfwcst2CPWFG3WBqFQnE4YPSk8Wb2T3gTGsu7Yfxb+QSuqSl4Mu+Bf2U1/JElTcA
vfR9oVvqTqPjxEZOSijVE5DbnVjc3SkEoZQl54quo4PitnpabOaExEJx/ot8Z56lJ/erk0kHVjTP
lpXQ9RjQI+m4ZxTjyKnicOoyWMMjfmlmS6NZ5xnG7+czgJTZFwvtzIZEsviBj9gVrRAX0fk7BbAw
JFbXr230CWjVUGbiS+3HP4omwserUsmR82AWSJvL3o54YJtkWW+BMIGoN98DUea3bMYWVqLewvAs
Bq675F8bH2Fsa3o1l1dxqpQ6+A7ZNHeluiR+4p6h8kf/h+ovsNhF5fiv50OGXFi6SDMOVZ4BEjdK
iveN4Ohiead6llkAfhn1Yjxcw61O4r3rYmzXb2EYsS/TslUELOku/EqE/5JKhJGtieXTGomBK++e
yDr3FJ/R+k2p1lgKWl35TGAS3cyoYEWP14qae2cg8fN1XwaBeM1zKi25D+S7fc6KigmvKKDc0zMP
Y79iqA15F8jvXPSKwFwzOHEEe4Dctv9LMdU6lYgzOKxu19P2kEBmfyW6lsFma29JX4nr5j6cuBhs
V6S27zzFdfSYSJAuaVm34V3LRPxDA233xlLsbjjlU2dUSTboAQhGaogDQwFSdaWYdU2qdtEv7gIW
Bcuvvt1TT7tuX1wM4p2cgpslM5QqgprRVZ3wYwdZONtjj/tvGRXv9eq+zNVq2x+Hzba/Z/mfKjBy
GMaifczXa8SGZlDKSDRkg3Cpn3BTqrxG3tIvsMg4YuzqAnYtkIEC+LPaXQdhK4T7UueSdT7OmARH
YbGxTg4c2WhO5Zu5SoQ2djDkuw6Xw3GX0VcKGuPpcfRyuoeu7SaHaVCHnzGajvJQ5oUx1f4kSUEi
RCdtUJOuoe27lgVLoKXZmP1CUVFIkloKDx7XZ2O7RqohEDwdYLvB4uZB+rcdFW1022m4DiwdYj51
K3zdesyyUljhaErEQv5EEYNAC5Rhwcjj6FsJbSeCz0c75qkxE1LkR9idE4/CxDE1SDzqXUAUWEMl
ZUXiUNgdXvwpO2hMvgLhega2E1kB6k1s5wHQjHTmtcbULpvSxZUnFKnk4LP6er25zT6D6ZqDMUVF
ThVxcUxX4+Tygf9XaedykKsSKOvHrBA0ss8woeEujiQmrh1DKmbwzVuniAWN5cw8t/McD9l6ih23
6wK6E+yPQCQohHOlTp0n/ufaJzZJFi0ROnlXHcnxB1ymehGtew9CwVR217amUhK1EfXAt+wqiRCB
JN6xtKOMOHUysQAceES5YbEjfDv0zwwwE3sORSfsxMhYP1IooCIUOWhOG9cgtDhznMsxGuFMu5F7
m1h7QrnN7vPIadh26pXwLpuLg7Dxkyy4Zlsh37AfjbGSiccbrZYvbhhmjZ+EK9254aeg1yZShr+S
IqTC4AXii9WrQjOWDfIqeEmasioxuZD25yhPkLpZVckWJxcWqM4CeE8OEVDkYadNuywUJVM8QUiL
bo18uu05jNirhFd6hBUupikp82Q5kU16NWZhfaAwguYdNoB3ghTtCSPBcNlODnYN3c+Jjyl+Pv1v
1AzsPWjNc250cufWzpKG2tXAVjupyns/SUv0sZIzwV1ZUa1c0Ph78H4BXGiwqBYe8prdeWV02AFC
F0VB/y8arc+ZTj1DfJAEvQ42St8b1gn2MPhC7inAntyuaJ8F/JaLtXt+gx9j5+/2w0RyqGNrdbTX
55OqpbrY33rTU0OJe5XvzJRfHjzII29iJfjqu88RMhQmt/N3jcTBjL+F2GDSAWkO2aW5p81TJzTr
s5gVFYUpmJtnPALGb6xusWwPvxzPoUQvX/7FzQ7KYtILK3XLyEgHHxS1ZwAitgXzsmB2ci1f5oql
yR2/wRvyWJGyBG3lQGG1e+D03cwofqa9MBHbuL3+7lUa9lp0oX1a/dmd81C0Qk1QYu8BTX4hEUXy
Mhj5EeLl/YuKRgquJlhuC3Gc66/1SX+d0QYchMXEogURTc+6WdbQ2tto21Rfwb6Ok8WGBqD+1Mfb
2NbsRe5sb0unjvtDOuvcj2Pk5FU1Y1PtZx8k8JrDqjWujpBzDxPa39B27yFCtslHVXoEl7m3i4AX
HEN7JiH24igp3wm1Oohc+IPOExLz1URVx60LlWLBtgG2HFvkEa7W+vYo4JuvmjkGTIlgpW2+/uHg
zSvYkvybNAQ6eaKs8QtjBuS23+ZQjVAYP8loNHnA2LTb68dx/80GyaXU5p2vpKvc+F1WN2aU0BUK
9Ei/hnD77ZsBeEl2ZIKBNPtyk1M4DPvbIudbyJsVObu12Xlakpyo8hfPoC9RI44bqkPcLVNjcKog
mJZRw29veakVt9UEYr/MMbEjOuS9QgCN8uCsidouz+DZfwDNKztzGCPWodvlppsNK32wQR4tJqpS
t0bIBEzsknWZsRdaKK0L1+w3t5Xc9PdfUq59lxZ3oLCkT5J7h2tBkGAL/w6IHj3jhj6AiH0Xa6Ze
dNiY+9qMgyTdBOG99qPcShWBaSi+eQlImCgTVr0+gFED5exq+EPvUC2GmJw9dcJniyZiV0tJPiT1
cJQIs5a+mLfFiwOOrPOVuiicXfncU4w+EWAAuCqR55ZBonSOqjwIdvWac4MsQsN3feLbcOIl7k8d
ddkWBTL5US6w+Mmb+Thz3uZAyCsX6PXJbgTaKajLvfazXh/b06NxVjOmmCg02K3s8kQPoiugIAFa
QKIzEeRPxOavpAMZyKVaBG1CgF3UfCac3sooEmsSYLIoTWen7vgMFgVZFbK6m/2Jf9IBzb7LSGy0
+Krh0U1R8Fj8wHtk9gNmS2Dftmiz6HpOTd6dNdvCDg64zW5JEo/1ddS9IaE0aPviiVkenLOEhQv5
zzR9UWLQHTGjFl7Q9fph1zuBvAN56+jF5fl8FGLMeiXT/NRE9Gz3CJBwlcNCsmIf8zD3v54lW1W4
UpYJqnYzQWFoIKTSaHVFtSvVUUuo19J46wUpI2CXKV7NoQ1ikH256232XeVss1elevxE4G/UneZp
QZV4e0Es+QX+18pjy47xyp5zCvdusrtBwAwTw3dkAM2BfM5GiZOVnuMz/j0FoRW9GdXKJIZiLtKI
HyLqN4oSOIOjnpoboHKO8jeuQRsL4KdrKOWWj9rfD9PIfAFfTYBP2cg7SRCAasCmiNjcVVpCRE7S
6RnSElR8kK+3nRblTQ6nyY3S0L5epivimmGkiOeTxAaoRKYb8Cc8PJExfOJcx1aNmLqD2f+Yj4cA
lwuYeK7O7DX+7eizSObOpdPYHRz4LpSgrTrTAbpFnCwOncUmLgM8LwuwpmvTL1dA3SoPNeO5mBQ8
QvWGjDK39bwRgozrJx+t8NCho1ru0cEnU6XaoGYPRnZdqpcCQLqcx/Vo/Rs3qMl6xsyBNRGfeeGt
BHL91G/BrZhEunjAr7tur78IBxFaTYUGyAP3wwpA4B5SPM7hWqDzuzTT0cZFPXiLlS0fLmxFY+Aw
4wwvPViUs7HQ/DF19nXLTBn7634PeEK9HqPzTaWKVP06bWjDlzy0yi2yklY2OIpN1eaSqy8iZ4iR
bG1vGdCGOxti4mSXGrNwlfKzJPE4Ki/UCiaJANLbw/jEMYPe5sDF1KH5tknRumylNWkHJd/WRfwB
ao8dE/HOwS0TavcTeXufnX36jpDg+zv9Ku4MHVluHyN6UTKYNlZNuNvKcjGBT3es1yu6QGqgKsHv
LvB5Hb5Z7mEHUSxBI0wCaycQu6Nt5kBzJxlDu5gAl/+KzUEnxzOZ6ufUIytBayCdQONXMGUzpzg3
0n2pyaU2quOcZMltUCZmBzHBPTb7NUTx0bEx8sMGjUgqUoa+nDJCKOzlbs1MdazBOyRupBemowSG
gYwdTHbAmFaYpd5hMP7DdkP7m9YmqDDSnOigb3e8rsIiG7dkOUVoiUUR6ZUzpJ9QSybxsRWl6bDh
7U7Okd7oJzdkkmPiB6Kiz15B+Cts7JoaRpIjWphw+j6s3yOQf4ds0y850BYIXIW9OmcfVHG70aLO
A4lNbUHUx+YddQ4GYTnQXX17+HsH458eRH8ewAp7jvY/FJf/ZpAdOkR8/nB9qG54Uh4Xhol9T+UW
CqoO5q8Q7EAI3qvDr/0ddpkp0zVdx2mPkqc88LP1QNenklyWeMmkC/mtwqlSKwaUMRHc13JhxwL4
oZtlLDtlQpNTBtg9JBGCvoQbLJwiBrW+W9f2KDwDk4AiAB/BmHCL+8wJH8pI+cvi64h6T/OFJDFi
SoRtd++XhRM7pXIa4tJ1kanc5p1Batu2MTqJwlZGeD70f+dJfu/ySL/gobl/1Vy6xm/EE/Xte9YM
qz7HYqHcV3g1aaIpxBpfhJv3L2kWfskgbpW4kA+66kbPQmxumUr7cgnTvrizKVmjQzrcSEKbpqEH
aVCgVdFrHy2lk0JtCOXKNFIKI4YGyvxV3Sod+Mcbz8CQN0D/6YiWPOl3y/CTzg8WvIVKGdxEd7i6
ol+J0TJ0XVmMDx3xrX1uXdiyAXaHJ6KLVdAPpZiHHLjFlDW9aTcLfTG9QEeWCPUlPeL6yTXYQoR+
7OvGWHh2uk4GG8S3Llz3EUpkPzXanaCBpcZEJucIK67lRSnNww14iFd5G++/UjJk8Ce+2lW2LBSd
xLCEWft5Wuw2kDYpqjkxUy4pSTD0BsR7Y8B4Lr4NlIutIKooInmJHQx3jm6gAnl+tD9MgvlEg8aN
AMmntypgkWIr3ro/UoFOso1DiqqFdOfZNJGYFuYl7ZJsbPWEX/I3cd2rMk2AqsBlLvgn8LgiOm0A
iXXZ8SjY4dBgW2SlUR0Mc4vv12uLHzVG4cMFLuDlJH0POZvDbaHWClGk36UOaPnSaoJr8Vt6M+WP
AS1abSoQZ5OuBx4HQQ7Wve0VpKndN4ht/FcYYSqEC93qk8Qx6iV2and+svd0Oasq7dNgyLHzvPmX
qCur4D1891o/ynkAvVqzR3Z1MVoHtSGnpWnTjw6o2hjIHZdnnC8Xhmvs17VL5GhAhr3Ol6Q0Ug1R
CW0DZZbw1UyifiiAl7S8rnmd/S0z9GQJNb+7ecP/Go25MJOdLwZVBKng/cvUhFePJMbtieA9I3nw
/rkLgAgnaefFuoW9ztpwO36Zm3BVeW3Ev+/2i5YBNgE/Bew7gv8o3tveIuzxHYPe8W9hjM2MjUGX
xFUdL34snhAE9SZFJYrrpBVbmAnhirbH9Q8DDJwY7k/DntgCTZToFZM/WpBe6IeW6NAUo0t4XeaF
W2zdf/GM+I3wRKhtfdXtZA5vOhMsrE+QK9G4aZIY/iLr+SqKWAmQQfAWNAdQL63JA6MTMxguLcxQ
l9nNL+cwExhYNswSPDAZgBKuMcsWxYpEm4YmHrJjBUI/V4rB3XvuZscFygPWGr60iHX2SUkBbZkn
M/OZSBnnWjWv+rPLMAxnvPxI6FgG9hxqz6sz0crJg9kZlfNML1b5rrSjmWgIFprKx0oX7nD1DPmm
dIrUG8Cu9B8qrA0xrMuw+itLunCSCi8TVh1GPYkDCnK2sqzVL98GgtDCk6X+9daOujtanNVkruGa
f+yxHUmX7cbBxaoGFoB/OQc0pNQ1MR9GntWugC7t9msPxn1WlfJT0j6pYkLmjdrr3fgyIxuOVkIR
WZguJR1eGdr5NWnaDRqdq/As9kViSYI9Y9wUQTHgOz/WQbqp2bug23H1H3IKjmjtGCupG4Jc5js9
Yi8wddkVU4d3wA9FpI3+lfwkV0Msn6gfYlj6AarScxyIkVyYNph+lhkF4qX7Fs0l8ziYY1SLscwN
JTViP2AL0D+R2wWUgGhTp1pCnZS4DzFib+Pr2TODq4+L5+av1kM8bE1Hk5dP9gSDu/iKa1n2vyV5
3xX/xpQ1C9TZjHn7AVuA7NhMwkk5zXbX6wkqxovATuR1XljWc1TIrlsl7l8cUivpKpjKTr95sYQ3
Tq+7bIJv7L7GcqbmDcgOedPUdY6HfewfCiccJInL4Ntf8INXM9Zl1V4y7Hnpyr07U2xrX55bqCvZ
1adPHvzgKiRym9DCG0Kb8y/zdvKmr1Z/fawwwJlXLpfl+2vd05hYLddV2H0+fYj28l6FfaH9vPCo
f+cLkrDgcG6IxVYoQ/tAX0jpK1lB53pDq+nkQensfQXfrN5ANS3Ikt7+xPS7q8EcrZ9FPOX4Gc/Z
sjKiM/kKDI1kgYoasQnGTM4pcr7ibtsURLwJCX5Nf95OCo21lM6tKZtbUtKUyvZdgNCB1FbDM0cD
x5YK0bAceVzu5oFW9kSeCd1cjxiMTPaJiEghjB1T2GII1RP1opitcdbrDuT4yi/Xjv+kmDDo7ych
HMKeT7P4IvDuqks9SBNw/w4mc6Ebe68glb4atEUxHFOHkynexTqQWie0n631rB8PLzoPeMp1cITi
pGtB+2wbLHz7U6Ia1ozEiONS/qZrfngWW/w8cZdGDinFwZTmA1KTt4O7hMQLhE5JIPRR/gCjO+Nd
Mp6lpexTkRYGUlzXMgZXL+Oa8LGylnfni5yWpBVY0iqgJLiqHrvsdQ/AUgov06ZopFV9paxVMimx
vYR/mIRkVi6gY5boTFwhLtNYC7eogd9UqAXJWXhW9oxkioivPN34CdFjs2E+3SbrktTKW1WpHaIK
yr+mKJXFSXXgilBSrC7CYcbY4Yle1XdwRkDn32SPJbXKtIaUOJdl2TyQbZg7WrS/f9ruGZBaU4G4
J+D+Ts/uWwB7gQaQ3ibDvnq3JWLpISC3js1R5DoOAw+1R4U4yCfxfAK+axs+YpeiprU9j66IeeGf
tea15yE4gaEqdXxmCFIC6SOyj6w0r9jMFCBaxxz4qthYUCqRsSV/y2hPP9hydm/w/482I0rXXBI/
nO3qONG0Zgg42f3vlSntgzT7aNrmf0WVqNNs+4ZHVCFwzcmTLodjdPJeODbxPdYaC8RiZC4NeiLP
3lwHXEnpjp7mQhVLpYono8igSCCk1neUJvV7ItQani4yhmkcu89xz85Q88Q83yXqx0uM9NC9ayNh
XF8yZw7WEdNyh6D65HwWh8U+y8nXPB71FwbOz5YN9rf4V5S2+uxW3LHP8L9UqY/tngpP6CJ+gf65
pIBM+bKxFuLt0WWknaQdEBTAp+ieAbpajHfeOicPbjfUgv39BD1GFkLaJZtCdfMuoqmUuai1DHRw
ktQDs++hsP85HKpgqsyl9L190eA3vVT3u4/fy+kFrzv8ql53k5Ki7UvJ0g75nfoTjL2dqBvZWsCx
bYCcIdC0aNFZpS2bOtZvgT8ilbq/ffQ6Va7C6maExs2lEaC1unODd6KGnngFfy7s896OS4il4Ote
ocqcdrvKoT6q8gyhs50Aq6gKjOSAvX7O4c69KaI/D8gHZrVogQBeIzkMd1QZXiCzFb79rZr2kCko
ktQVrsURQNWhpVIm8RKQmwBj9ipN8rFSCWQuU32L/0Msq37w15mCtjkWY6Vkb1KKFspPjsv3M07O
lFv401lo3YA9Lkuw1IRjQIhwCDZlkH1koz8VodJ5EsR4WIZBIIpiFO97JOofwmk0vwXQunYMJciA
DSOpNxx/l2SGlIED7mutAjSoLK+wXcnd0y+0lrlCrEg8d+dIIjI4krhiilvVRZrNRk5+F89baZCx
ZU0IkzlDl1zwXrReZCdIVITXT7iq8+wOXjE5bpf6yEJdwWBxv6LErzt/GXTUOUWCGVJ5IDhZUMF5
/tA3uATJlqEuFGVmKFZnJUWWWdEle5rPcq11K/ce8P+F/17nfdF1dU+LqaTEsO5zkA6aXIyD+Qqs
gopO7XZqBy9QcmS36gRifzQT30jlNUoxyKADVjHBLEUOKG+9VQsCf1OOrsVGdWRx0MyVZbTEvUKg
NFUL5opbd7xY38XMcQK2u2r6CTVFGVNOfsO6nld+9+eaaCdmWWUKkrKJpXT8EuYWSDs1nG8niEYO
y18OfPwQv5aVW9WIvdrFP1WM3mYYxKeRGGNyU/vJPXUEMKSKVaTJmebzB14BnTpige/nit6kS4A1
3K/X2nAXxA8iftmrSPxTTE6LgQJTTjGvxihDHA4lN64cXNIUU4RC/XMpIrbtNEK5FDTgj0Sih63s
lxBX00beKkItkneJKPlru2GdrRtNbamx9gtYYrl43xVpkzbzJSXQ7s+e8e0j8Z/YneEK/VDW4EW9
8fyzEts8p2yVSqHam563xFUgwQegjlpiU4da39QzUf5FUa1FqCHfT0XFux2qUAyyFwgcY6ywr0QS
J3Lx/3fGwRb8A0iXD9wfQSm9cY4QuMn59aNq8yKxPCAin3GhRsgc9oqTMhYctVWWcfvXUw2Dcnef
Tlcg9Mc3JgsmVC1o5MFTWEVMB9lfJdPFUIQ2EsGoGIX9XimMuzhjOfSti/GzRUv08HdgjqbPVF/M
HOOtbQjN1R+AHSI3bBRLVPsrMItzoiqX6oniHKIU55k9TzZGAyXXLTlHr9tcT7gRdQp8pSpkRlos
ZH8Y6TG01suJ1+7h8rDr4zJ4DokNm34lsBnkt/QKAvMJoVM1iZdANNu4GQXnhk2ZmyETIGtbpCHQ
/LG8veTkWKL7myOhd3PCV+Kous7lcYRGWkm4NENcXnkUwK9YPmHEito2rQrNMO37b5JvGO7yAsIN
7FhYbWncfWlzdQo46kK1Ko6bsUEaOJQQN9UEblLRbKDHYLQtRBvyqfU2hKiuojzT6oLBuAy1Fwxh
znC+hLw+Zo8RPB25b+mE23gshH6QPYLrA8a8LXnbH1gEza5lklafc/85z5eAiachnWYCaFn6IzH8
tOaYdu/QF+aW0nAxCVWC++ikfjGZ6NeoCUSJ+Ij4zckcgVTKRXfScYGer3BM43tBavX2+FLNBJCH
sT07evVg0MPBT5pyYKmlgUJEpghYlqwLiPRZi0S6tuLjUrFq6XBJ70E3PYdPykTMq82rkqdtIohQ
sfXFPFzmiTBYmbirEW6CHvKLsS/n70YncoSRkDy1vO50EMajSf8dCYVj4kTtiGPhP9X87NC5Sp9+
OwY74OZtfSJoZATgNF408H/RPewn9ZrVhDeEfnhroRa9l0ZGVbPARXDa5BSW/bL5CpK0y4QGcMWE
dDuirkPke7Xm4trnAwvnriLk8TNISKzgtdqzw0jsvOtNDhNwHK+VeR2ExMRHZqqF5dFUgbDN/+ah
hzf8407oo3UljLWtmm6UPJv8XkVjPYJdES1fdwavtAcnJGooUkNfOCGf/piFv8oZxBoJM87RFli/
SRDmfv25FGYDb37v9BMlmfOueMhwF191OJmjwW6gme/X8lzeN+p/rDsdez8/UWwdOEexTVCCgBdJ
Wy8tXywaWSlaLrb+RBVsh/7w3m7vK2UBQnMcVoDSKgO4FYKY7fxW5Au8G9pQT6E/Ct6Er2gGUnOv
iC0KLFH/CrvHRJpFd9WA5STSSXTlrcz5s3b5Fd+vYmGoMTxTHf5u854mCcJlE388jFrUr9kwaV9Q
nqPdWDydXlKKpLsx+gb8/wlEn5leMDQAeoGpRnphsIIO4I7/BNl7U8jHdI3XuC5iE6LPDo2QXHUF
VIzFpL6ZYmFOiyLe6vdV8aePiTm/48D8Dyci98l+LUqY8m/PCeVaErlSEs1flR54mshYg6ZY/lDZ
UlJNCVHkJLtkPI0kPDyNLek3Eww3+yK6wJ3WiMoOJASu824Ir2u1slNV/15McCGnRTxPuPdUcTx7
7lAdfui2WHkOJaMF+3lkUo7u8bzKzNB2wC/wvHnrRVuqaIEFmmfNEZMCHTQfXSnb6xeKZAf2cVIa
fRsI8RvGSexGYf6VpV3kkWbGqpg6t1hiXJL9fUcEDo1DsYnd/Q25antMQMjV3qMePoM/HQU+Zw9J
dG3w53tDxyW7bt8CT7sug7mNdwOVBCpM5s36Kb0TbWlAt8FDpHlVjv7G9diC+zi5B0gL6UXuk0zV
MhmKTrp3aPO9sPo3smiSxAIPuytkt9D6+dQ8aPGA968XXu6DYVqNGBFJuEAIOgeJ7UP9iGi0pG52
4kRLS6dHV4kkS5hw/r+5X4kpFiW/I+zLbVVvPr3LPHgdDCbENQD5LYBQVjBwlpBrO/hvwsUmgPb0
gEDVHyURuWlDDXvzhfTSIj3jajjSyU7SlzIH/I4/bwxMKDULIkWrNI2zuAVvXG3gWFO5khSIAx8y
Oa2M9VwyA4y4U0Wci0b2d/r8HpZX3dPeBMBhog6ASnQONHRG7Uf4IU9pTJRkh/ybTpxhVNKWP9zF
xJJRsT7MXD1TJAhYc3kg0M+x+zZwbvH6/jAgknTc3L+1ujapY/sxc02w3GgPYINMlHQ1mnrRBGhm
MPGQNIGH69DsqIu2UaXOQUSQDK5Zej2Uff1PM/RznZFspxHGK/G7EYKUeVyoDr/H+XxSdSvIhrRS
Plsy6h59HUB8gTONy2Tai1q/LWgUTL0xjLFr2yKQQUIXHvKzhX27uuulfCBal4YVpdNpCzJdjfWp
dZyD/P2ESMIofIblFXVRjRBeoVIXv76sT7MhqPZftMdLEa2C41v3McdkiFKvwd3Ct5xDmv4RZ/UB
Tm3J01DWWBf4z+Qjr8M4uOdvkRNoeyaHh6uNoJ6VC1GWiD30WrATfiabS7Ztp95Z15aQVslxfZfj
at4tgU+14yH+rUoeRjvt44AhOLDqar8Sr0ILz0tjyWKZkUCH4N+bOEwcVS0lPv0ff5vCwOMwnXw/
HlMUiwPeSW/HYJ3uixDjeokK4QmvghDIaspTR2gUZTN9iLDT3IiU3PE45LY+G8b6IP1faAko/5qk
BMVKJRRqQvands74o0rKtoKf7gXHDbnhOOY0yeLXESMVyicWGVBMA9KxsLD55kafOSc5pU7p0Zbl
k4iuHIaIkCtzwx9Jwr4MNZlvUebX8JsG7Fq5/7zEPRH8D9HejDa9tKFVp/6j654aj2jEpbNAP7PF
tjw00wkJGoqQ7E2qYzxtVGkiNlrJ03rXAJglrTltJ2CjTnacX3lQP66+q2fb5B58+xNDqAK9quqN
R0PerHEGFH5y4upz/fsPeN3eo8lgTcpHE8iFmQJ2w0GZiyBMoYfFl5j7yFQPKYw4YDUFUtH/o7WW
me2bSmDLuCxsTFaKGmokO4Ik6biZXfQFHbH0PZjKeiqw+NSHF9y5XDlfZyX69pcQN8I5bFW6AlrO
CE1J3hFsIAPkMNQEGiXG2zBG0+zlQUZvxJInqVDUuzM6IrAuXJMwn/Ii50lBcUmbXhdxFgyODB27
dZaKdP92xNkTvoTDdFeChDcl4fhYEMiQpuoKgvHHskzCHT5gwBL5oYsFtVmoBklI2ZwwNBBJHyzx
Pn2npwaekkTl+vuEpNa8zhJhbFYf7w7SFt7veLqNq8ifUJs52NM+NA3WWrg7PbPHs+r9xb8+ieRF
WtmMd4X64tFjhfD+2KrEB4oOpbozR5hRR+VD/EYvewyAtk/mHsutm3MHH2cBW1WiFCLykYuzJNNa
uxlTk8exF4olayU0ojCFBNu2ekS9V4GxBKx2wxAHP+DQTuSOMZ3c0pibPytTX65f1RQ9f8utOKJt
/G1jmrcgWsqavBpSgV1vjnZ9CjhT6abfilXlSIxGhAXrl7fMSGoL2VZbFgIKH9RctYoIDRhbcCzs
zJvZoMowC7DJDJetDYtHDyuJRqHOZfZ5kq1yh7CF0o4r0NGvVuIdDN5Hk/ryy7YLwp3jpzbLyWMw
zdnAPxppaqImiyb0fv4KIpvythUxfIH985qJ6rL1Sg4Y1DiHB9O6evg2WHaj0b/Oo5O9liTJVqfD
ZUP1t6NBHbQI5O+B3Z05InogSH2N/o+GXBt+I7v0zExs0flogVIglnxl/QBoWRXjP4SsSQbezWn1
c9D4//XBXCfQeqk3Av62HlujmS3DICykXeF3QBXM/yG24ireeqZdT8vEYbzbOEHcrjGc8Ej5kG5L
hcVyyzB8zDVnUnWXYKvHxzwg8A3pHdJfiFjhM5CfgyxTyMVFidF1rdnCv1apVuxdBvqBIthLN/nB
z9OK6pmJRFwsw6u5BiHnF0AGdangwhUop8vtzZyubl9T2L9awdXHDOfXO59uSWk+oBYEam5huLLu
cQwJVqSOv69ZbeXW6StcKoh6l0A6w4Yi/mYFY3xhZzvJJlxkElY98QeCqrPxYse625ygoo5PA+jj
s4ElNssDZ30/UChKdDbpX2mmB+treM8gbow6oVqv71juv9z16mBBr/m0AbDLAgqWD2+JVFuR9XAy
oqWe/dU/Wn374lLyqXpQOOftrj5W8CI/uGji0yFX355rMZhk7g5ggn0gHETuGXUr9xVie7kNE0MA
TIGZIomAGCP1UanE4xF5YxXrttdlJfMDKqywBuRcI0VOr9AOKpl7G2Yx970552J5yaf0Q1i8A0W9
Ti2wqE9tskHDBPJLA5pac8bvhAjmA2obIa07RPIbTKl/CHkg8CqeBBKFj9sg7umjwsyLFe1QDIWa
fCyytWMy9H6qOmncvxEGhszD8tkdQ5Jpu300wFV1nJ+EODS2T/z9BeL3N7X6O+LvD4lNs8Lj6Dhf
aJRQVM/AqVHYIybVyu2LoxDe6YQdcKzq5SanPjHHgKTQJkssa5GHYndyyc/6l5z3blAF7IZGScd7
jyPUS3LerrUXRIjUDV4Wkdb5jk9vV7a3HiOtZlMPrW/yWyL1DCVUPq/MfKziT0V9GrChp4DNQLBG
9Rwt5ZjAxn99Qk6Pr/hgxquS71j7Hg28I4s5a764K6DpzCH86Xy4Prveo+TegFF9L4nOClTV6TU/
ZfZpKMy9uJ8vXIAczNdkNBIEMSoiZokePffdGBLgO2pcbEYzIodkUIMePDLqi3uHIxtS/U3ImKvt
bGaOXkwS5NwvJCLeUd1WFP1uK2MqkX9Jk5W0I4c+wNGONeHun357/3ZXS54IgANfgMNWZ4PSdrWQ
vxIXaerYTh97xYAXJ0P2BQqiHzfmMjHW7mYeBGTm32pgDcDmJJSPuk3kYKnVQdMtoSk07CfP/COO
QOskJpNRrFWwCpit0x4S4bMROgMGXGPolKKc49D6F56Y/2hs7a9roQcPvXOrKyYb5sljENFaHsre
tKN68J/oIPer+JZG3tPNHRr5tU7NZgTuU4u0SA9e6AIw4y7cQ1fwXuADVzOOVeJNhqZRXyaVL8tS
U2oWbLfHd2JPZYEK6tbgpcInUpys3bMFFl1hI2L9b6pwya0bxam1g9phSIxM/5naTEwdc1+1ahHi
fopX8A+85JeEusOvq0ySbuBDHas0ndBnVOkj9gK1AdLxaXBOY8bilfzieF8x0M5TwR3wN7tUbs8f
up4/I8/Mj+i7G8KpEe6v4rTuWxM0qODs64alaDWiKfwYirMSefAYu8pD+m3g1Cme9URvlQ2TVej8
ibQzx/7vCaZw/mFadTG3N0nRV5RgGFd6gq/nF0w6js3UTVbc2+Dfhmbdz7wHiQ1jTFf2Y5TT2DOP
9vXcRLtBS+BAErej1eJxHljn1wPxVeNulrHDF55dhjcVx2fPVCNhpqNYV11/YI+h6Tx4gFze49N3
SJLPMbuRKRM3GY9/rv520K4JPd5xJ7ldST3lWaxhoMubUQNHhAYPcjywfsefq506/Mb4/BsL+hlm
SFvv3fvw88og+Fi25/B9EqVmyrLTAGLEm2qbcx3shH9XOFvrvXBtAHzmuIj9gCvrDTLMH7QY2z/e
+kQ26RJDGYA83+yeuXQdIhURQHUwdcL1AJAFjRTD5NP5NAfE/NIm8R+yQTaleq7SE3XA+QdBFShI
vNjG9M+8/HgkbhGcqy2uet55/Xu7Iy1GxzK5ITByFTvS0Cs5M53mik37fF7f8sDzUA4R4WY4nB1z
tpw9w4KBHL6nRXZw1e93mDx3DnQsT900vVSDthpZFCd0ri4ge6wGhGts38FdD992V2xmpcs3GbKb
6yjXFKxYyKPbxM20MwKJRc2uLgRFs9mvTJLXDDCU2bhOxjl8eq3XiDybsJDdVw7D+oeo03/DK2A6
VCFe75UURRG8Pz6BM0Df0r4i5q7S7Bc1jbcRHJk6dRaMImQVzAQNC+PEwTAbZ6/JOEqbH6zZQv3Z
Zg2sEusRpGP7r/6t47GDGawjwDIzrGON6Zf2mFzc8ALn35lVQzcJHt6/2lbvI7njpH9MQXtDgo5l
mVUXkrx0YULstaHfaJC5OJHG+YkRL2dcWfx4HW3gKXuyUlfMkiGUj2IibwpYTm+hupUhJPTGuTlE
5zNbxcTaDGGRL0iAFx7TYWeRqNPwzg+5aNBEEVQt31mtSFn1BwjP3dRTwVYSizcGT27GvKPrPUSG
4RKUN86QJ9KqNqQ3gSG8H1Q6WofTQIga08F3Cq9+eEEbU8lhrIll4O6+HsoAsv0w9v33XEWNzQQI
41bFsy36rBZ+Hk9hObkGudwcQqAhQmmSfvfoYFkrnyx0+YuR0eAYa980X0cEo98qmlShZiHr+KEY
vLTotr4kymPi21Zlq/mv6LmAraDnOmlclPBsxWIPVVdsiL0zDIOcQvTN3baFy1lTncdFREbS7Ujt
6a5xDZ08Pj+aUYJM5YiYfIq63oUO3uainQ8UyLCoFXwrINLV0ryL7HVL1835Y6sXblRjRpSJv0tf
Jne6bZRHyM2qJcBAkV+2B1OCkjB9hcVi58Y/YmmAdASS34M7jZ6bJ51h5fCXjv1TxpAM0if/DQWW
DVsyzhpoXtjTr1CLAOFR0VJgemyvgYjuXHCaOsP1rIHgpEzfKJJT2wqV1u7cfuyunOm1V17aBpHY
ya6p11jbA7xodCtRQvsCfstJ20xpZ6sTHfYOueyRA7OaGSJ8/6sKYclSua4Bh3Mw3MV8iZ6ARCbS
YrinHv+Sm4HNP28kmAJQrQ72vKic2+mV9DAZYA9DwoaI4nby7gbVvknaEmQXxdZZirpiVGNSn6Se
bCqNfnG7tBxI9iaEuAwDnf2Sou6ue2O+Ep0k/kLty7h4nQ9/nZd/Izeez+N+2qoXhE7t1MILrqFy
yJbltOjqMi1WTwUrudFhTyFh5tVA/BzqxXE5f8Ku7d3bbwckNlthQTR88oKNUZqbTsuq2ijbsleu
5TQeBim9VfwRMmJxBXv4A/St7ZGtcnZlVJCq/KWqL3SD6/jV2MkJyVXd2P0E67x57PYn5zIDy9Gj
gWz0ytg7T+rOkFfgamuIV4eARp3QdJXuHcee12AVY1mLs+HgOfGWqqTeWQiGsl15de8clOxbbhS/
lzGsFf9AtiqM2M4f+XSMDc58si+KNLJrnPCaWdny87KrauQd1eI6YZTxYhn03bEtn6rjMlzXiJbm
Z897dOLBctu47o7OLdAhslAdKSCof6fvDDnR8zZhOb2pzycvWByDLLwWV9fRaxkAUOy2lhhKoQmA
zOPgPJr1ssQV80p6QcqEc8PkhUNZWBkh2xP1ifCN8pCWg5HOrtssgYAP76wnW4t+nJzFKgw2YG+n
wtXUw0f6Z0dzz+Ozk2SJ/BXsP3/+F4tyx7HfjwdOvFPXsR4JSAMYi8nvaaB14r7SrfN0Ro6tdGzJ
K5+Y48SHAKI6D3ACpgKNLwZ6g0jyVydNvW58rzGo21g22kVtB06+DJH2gzpDQj1OCCWBteAZB3jT
3nSiAC2sOZmWNGX9T7fLeOrjASsVVmjyT7XGBV/hFllQ6F9ldL8f+p/9ACthm+Pq/wNL4FWIuBx9
rJpaF1gR1JzPdmzq15XA/33zGm2krP+ADh0n7eA4w9ce3wtgKa5ac+pP2bWAAbuKXtXHws4frKfn
t3cIp61w2RnzF8QDVuqDdMHktx5UWwpiBDtgf4Z732X3CMCVJCAHGF7U2nv1dFIEbj5O0S3a0hlF
SWaXZJDuir/KIMqNyKE2Xf47zhq93142xspK09NAtWczgJqYe0rMXe2Rp93fd6Za8YUiCedc4ajT
CF/B1IyFV2qxC0GTnaryhAFKUmtQbqfpdGgmqDwmQBxxNtuyBT9THaeVH0IJ1EQmsn4+3dsWhLcq
PfB52U4PRS9kq6xaKIxqueSkBs/bMvon1XNdxBVIcM2nidPbUu0qvzsMeCZ3aCWgJFmwig50tyWc
FHemDKN/4M0ohssWMswOq+wb/C+n1pZpV296WAhBYY2vVrXgKFcPGsOTD5ssR3ETqyItZWWGgpDV
enkUK3eJOHoqNsAStaR5tpIHHtlOUrPFm7Ip3BCJeoKlVtoL27WyegrnESRw/QlZbMfNSCB3Ru0y
YTSzAgrfVAkr9EhBGuE0SNcn3CeqKEwL9+w6r3WDXo8MpwTINoXd8Zeftv+nfnLH0pc+S8DkAObR
07YkytJHOWGbPeZkGVC/W5LivJIl52I+lcUPTRXqRiAX1ELgwEMN5Q9quIFEWYbzQaHq198Ig6xH
/9CHvgIpgBGfQXuwvvEFtxt0fyvNDNebaXob8Cjh+dP65czOAJ9iAEYIJ/1tgUhk6v1/M6yeYv18
88bFbQ1OVu+qEeFpGHlW8OVO3jcZLvLOuUqpr+2na1KXKfEDK0PlmWO1Rnye92HUPonVpl5QJbvL
npAMJQDV15hqTtjFAQxOqQdHBnXqjgOS6AHQYc1W+z8FGhWgR9UAl8iPtJR0mb9soHTi/b/HeyfJ
Vy0jRxVJXDDLL3QMBYhvnH6YhIjYd5hmipn0Mj67VYQlrIUnNUykinvQDtJHESz/8BUY7fRg9h4+
pdNAW7dnMgOXyQP2bqIUv72vhpONH7UQKGRbECpZEQWmtzYlXoVugQPhUX72vmJ5hJo9bsrJuGxa
2kZ+n/A2D4WW70kU5GsreU6x7B2aZfTqCJNOKzLHMHV7jzTjETBIKx6hJ2uVeLyCH6haI2ZmmzFH
zZNpRWBnuttGz/ttLU/8SvB0OSnYtalUcZKRZKxOaTtclOHSihCoWtVivJvMFXqlLep2gcTPPQHz
lkqCTCukL343+CLU0uL+q8SQtvm8bQgSEovz4/86mUpkrFF33hVPhGrLet0OqGmvPJ8Hq9EGb0x3
sjCDL65QXGxH5Z0o2agW8z3sNdH+qM3V9tZaI+/6Hx7Z93nENOSLz+9tguOKY6GhefTRLtVzrIoY
NI948k+yUnZnCn3P3vGVEBujNEeWUskG6ZyQ6A1AfL1z49dDwaipIVjPZ9UPJN5R1gFUJEWThslx
Mi7YBq+pjgb6iXLotfdZq47s+PQoKd7/zMBRzFsKevkAYUm0StDVY8GxE0EHKCWg21vukyE1ycgU
65oC6C78aXfUU6llY3s0GysT17WDWrvjbetFtuoPczD3vr6q4efRpgGgjekXNYJ8WieefJkUcWZa
/PPa4fPddtdzwReCZEy+teO1wX7OmGBV2RiyFvDkpiaZoWJMlwjgSIBPnFAv2yRBKqCReuIVSwln
fGyRoFXf2GPAPwqZpBkjI48+kcV6W4s9MI6u1yxJvVgGJ7ZVmoLafCX5Kpn3njic0UWE2i/+L05b
/+i3ySP33VMld1AEXbCDCPu4Bhuv95BxmYPJfP3HvsmJQ2FEEqAuEXKmQWWQZfj2B/v1MW8Rcm4Y
NZHGp91b87wx2GbO+WusFjwdWl7AWjSyo/W+i4bFcK86l+P+KloOBY3OG3B/DBJpfGR+aD34Fm5H
FnQdNlRiLUIeGafcQMxOr/TsHPT6q47+QjRIww+KfFUru6lz8OfHVbLklvpBKT1yP4C7JxvxXWjs
LAfQVOXm9S+o8UezxpkLIpfikDksAGw1o1SUKdXkD1XCXCtNzcthuy22bH4q80nNu+toENZrzvJi
TcCu9/eukxhZUoXJK2wCFI1OTyZpZZeszZIe+iN5fHPu5dn8M2G3mHaL1ojfHfF06eFkVy3gtKGE
sTskYE+bMYyDwkf48ZjHHGGXv+ShKYHt+eevoIL6cm3xiFuRpIGP/8EIE7nS7iig8e82PfueeRgl
ZWmoS6AzHuAbmyQK3a17Jdiw0zSH4L/l4q8X9biALEzIx9bV17tezsC07ISviNau6jbQjEVPo1JB
RDzSwO88KNGe/n2zuxbWU/+RVG5MTFcFaGOh58LmE8gFTQoH9YXHz/6DwAq81J6J51BqxKyDzGpo
/L4X2hopY00flyIZW7LPaXwp2SFS7618WhV4lHOdpr4v/uvg5vNzigL2rF5nAuKWNVbJCJJOVAsp
u32Q48EXV45YXtpZOU/2vJy9qoNJaRKnEdLhoHRP50mzJHk0m35Huw1iTi4mal1yJfWHFphbjTpH
hn7G0rkuV3BB2hMy232AaU/XHFpa3EU409TE28hJhyy2DgPZ22fDU3kjZqvM7Kt1sFWyxdgrF9Rj
YhbBIAPgPtlMtCaD2CJSSabbNlg5G/IvW04KCXJcR0JdEXMLcOvvxlCIM1Xh7ODDKIqB9A0NJLpv
B0FOwY0gBpzO8fL2E/fJN81q7XuLVcuLDVGCfgcd31UuGUgSlB7LHfrAACSIFe6umrAvXM19JsHO
fbtGMcRk2JD45sbThLTwHYGTkd/nxD/CWfbPD6cFhqV4ovIrmLtLRaNaPO+qaxssbZ3r+wgAOhu6
c/qpo7wnB8vPKmhPLuf9PhrIKQCqSqMMWOtuUI2GsCanTwkwR1SXXqm7jfq9X9vzYaXaHsXuSL45
weAG59V/bzvNQIGSO5awVXgQFPgQOgCwmR1FrGmhWWMxYoejjLLDWiSw3U4mx59hgmnW64PmsMLA
4UgpebRzFRDZQMmKEsdewlCahWbxcs5clEDP9uwVElVaUXqhW4fBnqRZsWmL+GPyxpMmAj/V2Ssx
RpLUxpAjtqq7iiHXYNmdQO5ldk2HMePqZIAqYKQJqgMt+kaiYhNonWaGvCKLzOJsfzvWKFLCuOHl
uX4003qZaenLkBlHg0g5f2uduQZl5SdTSzoAXpt0huXq4fh/isiFZSsawRwHgBQSBS5fTaANw8gh
beHi+ne+IkqrC0hfbaXEEdD37nhHYWfGfJ+vz9ZK+F2SaDxVoWPg2y/skSWxTRCCW1MPDEnZjRFO
zbSdjlTxHDQTI2wbxBb6Agb/Eyspfbd9J2+lOOxZeDR4aDAa08LpUDHE1dhjJbwqSyEcaeoJF6A1
fmE6g8iexcX2nD2xImHM2QlnouBqF1MovX96k0bcEUmGqhg6CpV5uayLDIUJyz1dWt6OkfVcXFpf
CVwvzOrMXqNjAQSEpQWuwHgSoEZcYSgUv8Ahdo+FI8BNDBVRKuHc9QZ02oupmKIHdu5b+I/khpBT
n4Uc3hM1j7tEVQ8FS+XyGVOh9VOl8OX/soxVrc2LmW8GInEojiOye0hjHzke2hRx9u1+ktxWWCnu
L7Lcr0OZfHT4pRQLkw265IaXkKd9OPCL3SNpXMH1kOrdI0nqo4Wr/xP2/glWkouc3dN19OAnxL+n
tEVUm6xcARMwyPuWmi/lyrmxJqdzkVDjwdC5j21YOqCVJh0GCPqRoKmLlywMe4sSk8Mf15JJKSBQ
3X8eD6qNJSbs+lpUaYuwkpt3kje5Jb4uXKDYjrYisT0Y4Bq3S2PadkRQv3w4+EgYtn2I28vXHSUK
ivdxT81zTi13fnN3gJiL+AkZQeKC/olMGp5W+ATDezBQ6ns5JQtN0t5SucsZJDcPH5lqHqUgVlji
uAuHKBsRtQ7Heq8SaC/0TvT+f31E1F4muE9q54FYe/2dfiGelflGmh4TBZ1qIl8w98H5jQOkg5QA
FbqO2YbhtBXKB8YWwwcW4kuftYwKsQeE2GIxFD8KW4JiVn2Scuaf0psBfLiy/ZZTTdT4Jp1aOsPZ
13TtaO2YxJyMr0Wx2YAKVxwpEVdtbtBDw6Dm4HUe3a+v+rjtVgu8mSl+V0PawM38oRfpaPkgj266
64UHmrk9ilHq/fl/acOwbf3/o1rrVtQ+tiTRisIEH0BzstaCdwWnisz+Yd6TMeg8atJtM4/9sioX
84JLiSgejthhJn0A1Hq7Jfp6EYZq9yNS+99C42GILixIEQu8up6FQ64j3sQulwpOgUDaFiUj6Nw6
lk0r5limQS39fIpegqHA88TL5ARI0CfNPwALFPLqEm8JF6QM9U4aAyx/5XGhEBKDl8XN6qKllRl+
LdePmQQgtZYuoe5pN04nYWtMB5VEG/OQ92HWYad0nFSUOI57uTCielYIRl+WGlwQg0JkqkoFJKEy
RM/dlIJd/PAY2YNDAibZ78HW8iGcNhvDPDcZwHdX9z1DVxpg6we297X2H3S+FubKpt6gzI6ddEg1
jrqpt+h2j1FbLhScyYCzIvUSEk8HecFju6tuNwc/WOC1T3k2CYQiebcko2eLidylgqgYSEgXGyxJ
qBH07clyJVedwy6LhbtL/FuTt4xz3fX/s/JRxMKZIaye+W+j4dP2z0s7cIZIR/n+91Ahat0EvOJ5
bcYU3OlLJC8Jdyc+g85P8C0gUS6SmjC4oFNG2Nsv3Jd3Z0bwrjj7uH6h2tTssCpXR9lUnhxwM+2Y
uKm7jXnaM1wnvGusZfKPRmfrHFOtNg7yT1mujyo+r9luBV/0Fw3CYa0kX9gsO3oIKKRoEis89tiY
mkj69Fx0Rm2QCHN1V7zVOZ2Euus6qniBi2Y/GcNGG6kowQ5dNtfufQ12AgnGMr6gTFVeI0ug12hH
XNLGUoe7KqENQfVF6nT3iBJaLd8EDYzc/17kxIlWr4u2Nu4TurSpdt+FAS/YkJ/yHHGFiwR5Okj1
vcGDbhUl0xIdKMde1ZIbCJJs9BCCdPxc21IDMJvOqktsXc608de+aipPintD9QWNnWYsIP1JkI1f
qOcxpFQhJZQ91djr/TGdwkJPJj3S7/FX5ISKBTaC2AcuQDWurpRBUAw88mQPK7vgeWY5vD78Ocnq
DL37HA4oMg2vC3u3h5qEgbs9MOwkk0zckST610rHvar/w6XC1YfOioG5+SaHlz2rrmQRoPnpK+uo
7CyN8UhxpCTa/AEKEL9MUDP0Cn0vur08lmLD5uCHltBRC8geIAzZKqmuWKbhDtRSpE3zpfZnHYQW
cV4GwqUnkAK7OB6zA4UbctIXoA/0aoZuBjkRs693bo4BXJudu7YKRDVf2sYJaaJmcs1PIAoeXjnu
f7yS7IT2VgL/mu4A9kRxMtpA26RSfyOq9HgEIoAR754XwxqCMuATSwiSCpbTb9oppI7QSrpvJs4m
ttZEFzW2+1umVDCpl8yldaIQtmTSCGEaFqFQZoIFc0GCljKlUSvYcZc/k4zjLeYOdRdO8As+rIcm
BfievWJhxIevBEMmVts7J78faXtYUQqlsOgjmUpBID/ZDNURWbRTP37BNgAb1B/NJkUYBW40ATDC
S+SZK6/XEOelZlbukMQ+SWfpxAvd3DOcuY2mDVYeStscsoWKuzr4rfIW//fAxMcvupTV1W2PNMUf
ndoMrx7zdObabJa964a/cZBfMtf/YciKS25uh7KmJwpupmvqTZcH9jybIROmR3ElQRTqMYrHikfK
XwS/o3eT1FExLZI94qR5/2F/SAZ1fr2HXhlDA2exDZ9vKUpliXyLDcHoVCSwRNZZUYy9mSeEUKju
4Qb/oDU+YHKU52hgOo6BX7d/h07/rXRwQfWzljajzZeQFF4D7oDeIn4NmGoxnfL14eoBX1TZKQWw
oBfkiYr7zYswmwFWH0EJei2zOx6KTgHDNOI/AWIFcysfNl9P/XxndvOnJ5FBvLwMqdQ5QG+ZUBnK
wXCJTyNL/FsAZiFAVFNsAK1q36CgF2fhNego5TtzoZQUpPKMkjyQvUi5nGSrn/OpIPll/GU2w8My
1FbX1sNbhjNtbuxRB1Nz03mGaL2Es9WesK2ob+5Vbya7I34iGW+4+1fPTlWrOpcdJzAwW6Ob4oBQ
xmSP6AxtmDIbj00PaydSRR7DEm4q5oLlc2x4OFMWFDO9B081q4m9LinPTvWoDvOh7l/tXQrxFsGp
8SbJ0n71eMYCXoFWsf+aFFkHvhxTqSiWM0P1Ly36a9Zk6OxfR+6pgxC5u/fXfgQedu2+2aZdDz8L
HHHWDx7S8YQYB56z5FrkY7JgK8Gak7QLikqtBtraFW1W4yAdwrESXB/HDUmLpidMijBm1LA2cNLp
3IY4rPfOvyRFom4pMYzThzflbJfZm9SBIainHnWUBD2T7z+uAPyKYoU9kkTE/moAhtCbTKygC2j1
obf8xVvn9WgGZAm3za+xGXBY3ET7SbztVaq1tZRgDwPImcjcFgM53p2GEWCjH1UwvEoTUVjt9gid
b0ijk8c1gTHZTpP7d+AyjcbAMaFYG8isTijguRbFFoWAeCPzvLh3ilfoIggZcqJawTLsS6K3fmiK
CbGJoTOO3MoE41oZXy+cNo2d6sMveTDJq2qAjEOGwpuFIhBQ6+nFZubVdONBlHqkxqDRpyy7lOS5
2xZybEsIot14/bqPMqZNboQA1HIIaZTu866E30L9KWMZJ10siYVa7kTlr5udIM6niaaBzrUzQiBx
E9MJiEnoHM6f6GLa4SVwk/SdBWkroH2JTo5quN3h+b1KsSOEW6/VhIp9r1Ly27B//RPkX8P3zr9M
DxIG4rGqnN611sKs+n+akz40SNkV6+lS2QntHgiImC/0b0gvlo/L57XevGeevn5Zlm90n1uAe+pZ
Ax1PHDZjzqvUphalVn4L0usb7nbW7TUzzpkTcaefm+cx1V7SNXhT3hUQbvd9ZmM+kCNNF6P6vLjs
tACv7H0dbS5EEvXnwpY5fpANJ6HhCppqRZv4hiI9VuMYtXoDw/Q9Fsi+7GTuGOen3epX3MBXCLh8
GKP5Kdd4U7iKGzgzQHH5qi6BM2m49EM7CpUfg9Z/oAtS0fhXJkrDySrbvzu6YmcbhyeLqnPlLexS
/vFRj+udzS7zg9jjAvnvBUzQaMoO8LVURUbUaNGVgdAgLsSYOCwWGRZNvkAQbx7vRMMxuhmVaywB
TbvhrctjbfX5sNN1W4X2Ri8uVi8SyM6hBtvwVV/LCZ2XMPu1FfkTraWtQB9jrOxRApSn5fW3otR8
WzXtZlSviU4k9SOQt/j7j9OLAoPh/HUPtiRzK3bflZqFo1zCw7u0rmJ2E9s/E2Yd/XS66svO2nYS
flro5h/X0+7QiA8XaLe9QN0DmLnqJ/SSM8bU+Z/Ymy6buHvd9bx1eUMol5I6Ymxqu0/K1eM0jFXd
/e74E+A0lWjO5Nt1QmGOHfHoqY4UE/Ib+5K80MYRbmO8uTy7Uyzs7kTZ49DeDcj6aNrxKXkkRJs2
NizIS3BE/sA7qp3eezvTMIWPYpx6zR0p6aTAVGZV5FrWh2HUhbrC/uLdJETd19t6E7//flqXYlER
UGvLGzquOBWnitXhDSoWUE3pH5nunCI8tQrOOcDqa7J0JI+x5pRV8xHGYpwp/JvY0BHzhL0Bc7FT
hbwjuc4pszfRMwACbPRkNVE/FqBfgKaIXI8L6Po6uoJ/KIU3eRZzsQs4D+7jC8kBZsnl8pEPT16q
qDscO/g9XV9IQlkCTZ0JH8uQ+d1PZnzg18CGGlP1VvCPcbqVpeu+AxgQE9GoML8QuWJZjXwHBbfa
DjP+wltjuMCcw9aVGR7zqJIeTKIjChJzPOxvt9ww3zIkVCdOfWhehtI0eQ5kSD5wi19esMCMgzSi
9t7VTA+AX7exIdMNOTfdnvxTcLSri9TdpEH/94ej25ictEIeHl3LViY6HsmFBiNZEY49YRuomfMX
rTDE7prjlJusxFt1ZiwcAo7mtXdDyMgtTaRE+QvHmiuV/K48Fuy4Y7x/2DJgsQBxxfbGebTzjSNm
1UrYmIKxzymeNKbYle92nVX9XigRFydomIJiPxcH/XlW+jDPwrU0MWviAjZjsddJd+pD8/+ibpZT
TQcIQ1oIc0Gpn9sLcA6JEE+1vX95aQL+RdhD+jIYhmzTqRjcJ1sJdZJcn2rE1F0JRKERFJiEkFsh
h+utGo2lKlWaC3j/Ke0Q32HzzREBpNqPTEUExGnKbDI9KgsQYciGC1j3X6Pkr8mkGXoP+BwyJ1mR
oDcOKV64NxLFhtNiTfwQjNdtQ/PxLbSTAuUfutcn+WX1xEi43G4L1DlP8iFatl4kb8d8Vp/YLhgo
AHlcMVgAuk85+SiA2kngDdip0wi40RCioxtA5e8yac44Y0Z8pZzUY6zNKXmDRXxgT9f5dz1u5R3P
kzZVRt9wrTVAsHdgQUvU+Oo3LvSQCptF70BPunYYJj6bMYv6ZTuWbj0Vafd1Bn+Uo6/XU5wETGOP
ehLZjVrajqMgzQ8EpcI6pMU4uvG5Fey+Z5xnrjruRVEJuhlf5LvXcxbnA6khJs4IZseIcPy47m7c
3A3xuZ1HSYxKUZqCOz4poXiaE3igFh7pcCmbtUiA/F8iZPB/v2EIcLQZlrH/uolpoCKCAaA8DaYU
5kIjQPuxjh/+Xl7cKpj0U8jBoKu90lPDz8pOSYg+w0/mxhO1xmx+uCNmhGpxzHtRUw3K2a0/O0fQ
8kQz4Xr7CQXsd/3r4QdIo1e62wkVHKxvHuc6puZc7HeF6HVIM1lSGm/ZkX1RnKKBYy2lfcK3KzpI
+5BFOBbXCtFSqnwkPsxxkArATF8bJrfFC9v0mcqco2V9wdTBmZu1Bq/KpoLE/dhsdzBqgu1LdtaE
AhXhDO+vj3gsLaBCWNHxfE5aqsLry9C+vpvIzfds6YI4034r0DWYi9bMNeQ5+5YJIXlbRa3Pkr39
DQXOEoBWI9e9NtDEZZ9U1M4bkrFM66rGFb0KVj5UK+RL54xHu6eb1eB5VNSKq0NCwy9Lp+EN5m2n
useyAWGl/T55aOvb/TGw5Swm9YhG/YfyTR6RbOR3wyaIBQ9lIE3gj1wuMhxgyAU79SA/Apy7xZqv
BN5ydZ64g5i+lP/X2S9hE3+L3N2bFSzRVxGEmTxUuarHTg2irM2XTyizcFNdnny1SIH4srju8/9n
65crGWYxEpkzAR+pLjtKrrEuqtA3L286Q4lDZVlC4jsNPFs9Cq+GQNMFGN/a4fTqsIBdjGYOEMmf
cQqguG6+bCYfECu8cY2LQA5PZ8SRq8QJaZDvkQQRHW4/ESxmARMGLEXqIXsAbPXxGQsolANgpwo7
tsyq2Oo51giqwuYBRBuI+Z8t5jEwlucEE4mZsyKW9xPLQunF7nghifIfno0Bi0/i57fQKEXOao3N
jQn8IpV9WIkjyXb8BMSzu42e174cVjFnUs5S+z5FR4MSANX72OEfTZENIB02GfrBLenbBpoxTwuy
iz9a2upeTakl47vWjiQIe6DPakC8cf6kivUSVofXpZpr0YUCvrjOfXkT7vz8gmTj4hJtf0ORnkoP
ITxcOlyOH1K6fRZW1TKUFTDnireznoi0oz8d8raR4xWAZZXoujxvV2psaa1hw8/s/MBl+WpQye5Q
0OIvoFBT9aNg80ahiFpVrLa68OaoXO3SVIf5Vdm1sysx/BuOZopcw1ZY6x+uwZH8aWEcEG3kKdVi
LDpL9uAsgG0xt8l15gAwR/VEQRzaqQWmxwnVmpQrS2rm33rIXROrDGdUalzFci2AuOQBfgpmkww7
vKcS773DlsueknKJ9n2aWMndGIW9O4Jjus115pdVLd1HzFgw2afdf54WM0uOTJxZaLC5hGfX3PMO
H1x5qBlDRTuOb9J2rm40UKFy+0sJLF+XOLNE0ENi4oYmhdGgPG1Q6e70YKdfGLHfa0DN2MLsj3nD
Z3/30atI59Vk2VHk/Bripfyee5yY0T/4FialG6POYY62DgDMoXuHqvg/vYPeKu2AR/b5XOchNq+y
KHzH1eTKCfaQSPePmg1vFc171eMKF9Wj/SdbOKfseQDTaKq6OWf+CrvjmsbijoToTWMfuUT+Hpe1
07dWdiZCGL3YtCKx+qbTsGW60Ql+hRtOPJr+R7Uf7tKTsTQnEiFewnykWXBVM4qHz/bKS+uPpx9d
k0T87LZmiVlOqZ4AUuTcHidzJICJEZV9kBJ4rsZOh28ImQaxYJ0TYIMIN4gwCif62zVPBW/N5vEs
B04gVnN573cygz8hXhyWGfN6Ufa+EZ+iB0p0CddwAo6UA+1oDLnCH18UMGXGJw9O3l46ziFB/erQ
559cXhR89oBSjplm6f5eyCASClif3KS0ZP1QdamEnTf0xjEYWD7meKa/Pxlvptw4u2yz3biP2cFj
KHXtunkbuppdt81bb5xcqw/v9FScy1mTOYBXOpWZrLQNQciDKfVB0AVqVYs+Rr/Y9HKvrIHtj6Hv
lKkqyNlpR+a2jwtcEds1UYGH9xCwDSU0+j5OVg/5FNFURHaSeBhAlbxJh9relDISKwA/E6jSYpZS
xfQQSQL7uEyExj5HoP9PAVSVxf4mDV7fp3nfG9mK8DYEYXGXabEcRD39qSrHB5f8SCUjBz9JGEf+
d3ycICUjSeOh3d/nGobMkPkGwesdd2e7sKJQ2/DfDmqlWKZeJIOkzXWmZHP/C1wurae3i6w1hEcJ
h8OEjM6hyudTplsVlw84Jcowqwac0EThmzVxjN3btt4nhmrAC2g7FU988D4JyfxSMeFVElbMmGc0
mS00TPhL9tfSLz1x/xRVTSqtpe1qu74osKqrY2ZP0agiBPe+uMVRHyThO9AgWa//Z6oFEWkaEh5/
vlFHBJbU1GattldrdbM5qzaSK84chfKTq/knsorZPwFjnS+rui0pPNv7RSQbFCrk2ZVgNGs8xwQB
zOLFs0RHOdX4jxqvUS3w0+E+aPMlC09sxDFU9UfYKy/3r+ckgUD6fV1hcfjh4z/Wgf71bmL5d7Y1
63dYfGL/ayg0bn2//KZquXhoemqR0keO4Hl5amAnUNkRfOThBK025Pse+pRwtAhUu2kfI5zkK9wK
OlranhrBzvf0TnjTBwshIthizMpNlopt+f89793Ccson7mWba5ZHnbDZpT8bR7p5hHQTx8MhCIoD
g65uCAH5TWxFtYcx4+nTgBYS6lRN3BArroeHOpP4zfiUiF5jT1q8XCm3o6FbeFJQ9X0IywCU6fSe
mWM969hS9jqbPCyGOZHGcqd39uR8H8ZMUC4+Ew/gni8hqmnz6vw0QnmDak1CuXYhzWLXN8iT2dpd
NQkJ+7zArDdTGIx9uquywLVIKl7MssXXOQL9bZjxhaerv0yEolFVAlbispvoj8B9+YyGfQmqk8Al
OpZR+h/LdjQSLeHt7sw4rbhYPWY73tL1QRHtgPVDd9R9PgCy6UTaW0d+LDU7BujQGYnzr4V0JA9a
vlC/Tjzbi8g7kiv14TYrRMzPxpcSGr4F9wz7SUjM8O8gpxf/7lbAMzBB9VWW1QTnJOUaSHJ6mXx4
mkNNgh1qfdF4gJcZQMAatQyWYDCdOX0mohMBYc5RJyx6K41eJUmzZBuLiB5Vmm7MXqWtILYCxhz+
7wIqU++zTvbmCJvZYn5EXjZcpDQEDFg0YgicyfVMxK6KOd93odSSNMdJPVYtf9LGi7rTC9tFZEWS
D863j4tZ1Alfs4l0scgl+bXZq1GGvEfkteocFm6ZCZop/pmabEyqMrxf+LwnsQ3eAZXs7o9o0WXI
sPeHRnwhfo2fWca4IEqjLBNhiFJPke72cJPxZRnnAx2MwMvafuweI5A00x8GqDFxgvQbsNZnhVKQ
OBUfoUqMcJmtniIOCXZgKreLdwiYeAnESbWjXkWLRJX+3tpl1SiwwrzS+H1tF58gqeIXP5lh7kkM
plRBdlJ3oOQ/Ji8ktLhv3RsBMJFXpSBLGVscnCsFj9ZzcSJf/Yx8zdyzlLnTJ0Iij3OGBPv4Je8w
B2Ki3/pa7048TUNeo4wQdKIVs7csLGZBQPUq/JtKVOpMX8O1rewuvczcCwWYUv9WE+vR4VPCDlge
hWYUj43XSQEtipaw687ZfYrU+mtxNFZeEotsa0Zib1P9u+weXtjNUM3vHk1v+e4By3T4lu7x4/45
+so2MdChkWJW9UeQuck3zqXzCyDPNbabtsojzuOnM4a430a4MEfJ2289TXcvDxEDp3pfBRwlOPQf
0BYTpmGArYG2hWmwMRYsI8iqwrBGranidNqGmhMNeOWKhbGkmHr8u0G/XctXr2NJK6zOU0k+ZIpj
GyH1S3PYKC6UowW5nhASEBOIevp0TQwSweTEhZOGayeh3aeOlkFrJ8y9msqCPAesDjy+oaQ4z4sX
48IpX2gnKEtBXaR0ykvdyqPL5HXOOYx8STuuw1IKAhARsNLkx7t0Bj+JCNT1spzLxgv1xSKg3TNz
niQcYWxY8PODDsezl95Fe3rqoqvTYyYd305cmNbOuB4qUQjlumitOOP5BReb35/AgPFIN/2HU6IT
NACBVOw0+wJNsLz18/8xfGC+DCL2GAy52KlN9vq53/WtrwjXOP20f2j9FQjICdT7Yc9M4I0yisrs
vK2UFHZTgY0b3SdYyJFTB2J2KKux9aaquINkebSkvIKaahAKM2tbpkWtlCKonwHoyUNRyrd1P8S8
OoZqWfwCG0ZCo9mTgX1UMXnXc8sFdQxHXBPaVt5t3WdvxESUxzKPxLOzcCBlWCRpFTW1UEr+rlB8
AI5PgCidTBzfQSLRcvfEaR4EoYri/6FgEQ+vKlKt8NEFTYUdWvgDRjzAD0Nrz+nk5FOnmeC5vleB
KyxR8TfD4eBnuHfUgvT9UMlhvpPlN48CEbG6JnTWvCEj0+7VBhyZiXPvaBX0NTYYSSbQEK7GS6RY
eM1HMmidJYxd4hMIdTjB+5m1PE+5vnrg3Xa2IBz9fhonzxbNzb8k5Dq9g0wbbcJg3lSdqEZKlOEL
pt7TvAfiLSTEX57bpZRRVESLmIQl8sl3iMWbKwaC1NCRpum5uQH7X9RHaKK7J09h0n+Bv9S4hTT+
EcBYKN0XPseidui2m4pQs8mqFA5fqsJ2+u9v8iHF9UyE5X3csEezpA5HJ+6ZhlIAdpxXE44g33Tg
Iv/9KWp4VdrtE3lyLgDfI1iDsow0j4H+frxrVp1E5da4fW2XWYrOeZKtFQOoNjGCjkIPeYsAGKFF
pMUTwNrFDEuQliNCIurBe5jxoe4OU3IlXy9gxILG9KS7mPrnAljyNqrERYzNqnc7aaXt94Jd2ic+
bm3PU+G0GIlMasTVWdzoYzU27vyMP1Lh9WQDwHIEuz5ulbprDsrXjkXAIXpRINYN0FoW1Wwii9dl
74zYdGG8PZFO9Cu0qfGU6HZ8pcrG/pP+wUwRRxqrBViwmnJLbzgPWxbKZpCqbhsNQD9iYgQCyrir
xkkJzgD5CU4gFG72oVIAK5QU36usme+/tTOcGNXduh6/ZJ8qcSmISraHkj/BairIhAL4HW8iLe3v
f2NpaVRLz9GsR+Dpm/w3slYgYFXY/GFURxAH6kqFOfA6t9+/uRZJXJ0adJvJhphCOldenCeQHniD
kgLgM/E2Xz4oMIh79WK3ZXWGvHJWOI8wiwV7hi+/FVqJh8Ng/wDyayFLOZgKy1HQduzlSS6BuQPK
kWCf5hvS6S5lHAsg8PN5EfBhzABTSuT3PREcLkXwaL3KqQQiPHGIGJNW9m5kFexFLPR4MsE84AlE
iU4UiU4UCKfYkMVTGH5dWpiJU/NLobodDZ7C2OT5paJSB5N3lbFanKzZvB1GmSC8AHYymSOwRdRW
rJYBOWB5oNuThWHPyd4G8qNRtD5d70N2QRljvMVrHcUD4OvZG74Giuec5BbcbOzHVY26rcAs9fO5
vK9AjZZuYiENXVmviVMuwp0g/i+mjWxOKbFSukvdp9U0BMtmkD/rDWTMpKbB9hVxbHuJCYs6MKyp
x761K1Qry1hadYNIzqUgTgu5Sco591c0VyrcxQmIvRNiaIwWFg4QIl57jpo7qsNe80vUzAuT5UvZ
OR1hoPJwsgem7YhJRkuqlY4G5bjdi5G36lLt9xlzKAoBia1Bw/+4m8FBWuwSjMIGK5jyxg8heEKI
72ji/DZ0DvL6dhoLnW1hqb2/MqHdKvqGh5A9TJJ5jO0wreOKxj2W1hHEtawmIReZWtt9Srg+MK2l
35V86IDZIiY1Zkp59IKHL9CCQMInKiO5xGhD0jP8Q4FTxvb/ey2QDYf7QZ9uSMNsH6a5PDPioD6Z
NqaIR2746PDQUoVWFhRLdYc5kfYGjTnWsWXWdzLw5MT8biO7n20AjVOyf/hepruSglDU0LrZmM4x
jQ7+29M4fKFfb1u7+VsWO63VjAgTV3ms/h34yVwbyLhfq5vGsJUeWReFDYqsSZaw4Il5yBpjvKOa
wXIbSDy+1SIL2yBhODI5tptsjNru33H0j31NalOZGOrywwXq/O4jMHrNeKIKVomNWtxiEN04i6So
w6mPqTN5YXi41nKVlY+25GRJx/HMtX/yjSgQAH3zFoV8ZtyvJklK9BheJ0hxmYM7lmFTFEm0Ywft
iBu+cfcFuG+XIJikM8Q772SmLXGKA718+StS8h9OxF0FvGrmI2CzvpiGPj6tjEioM6eKso7hwEqK
UULWqgUe03gSF9VnoIHahXoaQvrwjlYRq4A56I1bEv0cuXrTSqxXk9PrQ9FJyakrmc0FGZHJGWY3
x5lU1L5l6L8KwfeskRcXfuxlxc3B+08CKMWZ9lHLW7060aE0OndOKGrrTcn+jOYMvmjSV6XjjEpU
fmUDJMJWfsntj+KlIjibhehY2POhMe7G0Djpp1f+hREY5nPVSKdMggxNlePH5rcEcs8Njf+wwdA+
DjfGzY919Hv1l3JmvkHPASOjR5Ts1tLCP1mJ1z/x7BUB341XcWB/2hlWDlKwOjT6pg5C1UgswUCi
SqDgXzkHdyg0w0hJtC8PdvKJOEJQgIYERXNEYMULMY1dAGLxFXcohxO8koq/IWbz0NORPEffQNZS
NqUtGrwISBC85YL0jLgHoNwaXflirt9TtzhXsLOD56qxmXBmwogg07LbZv9gLSfTTRPoLEmehRgE
1TtObnwfmF/3drvABc+fUkuZLIs/cu33pFsjr1ViLYR9noLlJFNzcLTltdrb32ggkp0bgygDLu3B
5wif0O4HXycfKpgFCa/bCqIA6LsBvyhJOZXGxKuf5yiIP4lTeiEOVMOOfSOWecSwJggGKkryFfn6
jeK7f+Cx8Cuv8FnJMoJ5o5d9xp7fCqu/tASTzA66Q3YrAgxyIcP9pHmWbJNSsP3QvpSmlSoTb1Kt
xbICeHGwInMg4FPDXEm0dy9uffEpugBdc4MbkLJj1dqpAx+8rURJe5wNcKdvLaC6AA4S/rBu/pP+
mNrh5mL68SWLOM+Sm2vwYph/BjdNjsL0kvaUO4zonWOpi9BMexpXHzSSaHYMDH2UF5jlg+TyOxDX
2vl6biUX/y345S4/97cMuqah1j9WNmmLFSNvLbQlOQZlmLrwQvSDnjAmC3nUTkEUSUyFT3JZoND1
DgeTJTQHVv4GKHO0fCoDzcPuJgPVtcgG+RfE+WmAphlKLh2i0vlCejdPkDqZNkpFEEQAq+5VKGN0
BpVQsyy4yU6QIqPt7hi8mrfp1ED59KlHa73N+KlNCW9a1WfLrnoS+HPHQ9aNR6CLFh5ata36xfGH
mguxcuveeQlpsR/UFJGYp2ZJ/PIqHpVlqoXSFOFQIVMeofLfw8W654sjSOavgppMiP9q1YRLm+Dm
QVX2Y8RgtUy+7IQJAYb07yrR6/7qYkhwIrhZH8Qnqc8GWbMimJlHghrpZZiqyQAVvrDp2TIoLjY4
AHUXrRRKR46ivnf7UTy7BiRfKVV5TemjzGxozn2iTKuni9mDl85YZRFZAJ0etY2k/iTW8dbCTO0L
AbIpnrVMJ0HsDDDuMDj0F/HGrqvLlb9WwarGZuCP6CWKVwfVoSu2fnVcD1/u7+uzfTUTuxTN/HSc
I4kbcWjRPVsMP6TdNWxU7aFd0Xutfq2fMS2lAPNLSxMUDpWM5HJuacL8vcn9CBIxuz072bKcGr33
xDV5a9KB1hFD5m8lvuJKsh160ow9Fe0PwHNz1gnOwrUZwlm1rVFDad9F70ydTDfF+KsjBDV5yhA3
2t0v5YDuTXNkSpEzUsHxZWjDcUUudrAnYA2yrqhdXtiV2AIXR1il9DlJCtn1rat+LjAM9+MEWJHa
Nues9GFgxuXkg3ZUjaeDz7/s+SEHKVTd6Had4aQazfrQ3NK3out3U0I+tLIQVP5AUrH4iOzlLaS3
w7j88H+rMTqXzexO91CPB8oVxD651C/HO/yGefTSj76mlUnTb1epnSoJa7QLn4qc+xKkICfbuto8
IOVhFY6SSnYqZA2ohgH4hkExc5g/jr5ouCj7AcfscnGI9IJoEI7yBhKlCUJYWondYJcvLVE2E6ak
X8JHBWWA5OboPq5ao9xAk6GYIsk27VcUNbONG/iLU8XXg2eKbGTVOu+m/BpjFX8tmixic3hPvqE5
Ot17nveaFrxDTcDMVyICAFrR2iq4BZR28IAsllST+nczBmiE0zu++38V4/gD+oZyJpCKOUgFOBk5
RZ/iRTOH0EOcH+sL5k3YOdxqs6V5FM+P7J9MwNE5Gzo7y30LLZ8gr+Zwh9XovOoZXqG8D7irj7y+
rBjq/XnhiDoygTYgUdBZ4OFPUopuAu8hGhsc+fNsqmM+ke1WpHtp61XLNsYYjmAl4LTRyiuc2dmC
pyLGTngZnhdcu1P4Oori4n6tsEA7laSHRfsA8WLxKfYk1/xYoZMyHVGGd9FcMSIgjT3jlBF7pwyr
hUlj/sDqH5z4Z+OmvofIZM3m7gkO6QoBeQGDlFIG4vE4h82dVu8xTJUk+WZBnsPXgu6h3OJ7nYZD
8WPfCwDkx+J0I0qjvDYIGFwyjPl7SU5QI9iuYbvphqTIioKtrMJwUkvaIrx4ZRcKOOQtyY9BCVdB
9K7u8XYgIa0+eoerzcaVeFJy/DTmKDD1KuUWoKjSOjJWtQKfUKmk8MlPXUXrvtDXkliZgnIVLt9P
3QmEOfco9/0ZDj42kLAoPjOZ5FYC9ko9mjyOaIphcqKb9cHMRNOeWULE92R4QLe10Tiz5UMzIa7o
WYUWsLrsi6qZIa0uRX/jVuGGXG4WftqSVB/FQaZMSyz+hmu/Y/gk+Ai4yMKKPviddRnjD1i74rx/
NlCiVcQ7kfStCK9AsqqHDzaj1DVrR9RywUjKfLRJIV5WlTTIxb83cgdYJwi5nIUc0QjxOqc8rkaN
gNXuFecoGV4XOLVslCLLAmP+8DVYGcBslayMHuXduXJt+Jca7nIDUW4AO/PkSiQlnuf00HzlE2VR
QoqnIPZ3PMw2JkDqihqRG/AKQ48KqYl1fwsUEcLOdQayM++9ljERDYTuZRC1zcyww52+3wxqFYqQ
69wGYZus4TycyqCTeuCVFQGPr9DW4akP2i4R/lPVfUw9EeDdhhVf2IMBHEHoCTKfyiVLLftbhyhM
Jpfzyp7cZNvNtuRfIG5dQzUeQOGLGYNv4yz0d2sY0HYHbOEm775kcdGLtmW8Q3HXJzM9ixWNxFYa
VXh5QQDvMAKH81zBJKbhw1Le/OvQr/Dc9dJtDqZEDhQnZxG5MGGl8NHNwGpEuCF8NhdcWCGAYIXA
/ukZW+RWA0oax8JLF1esKWnx71wTstBFMvFgAt9N2A0JMUeIg5YpJoSx/lUkdjsdjaG57Obk5d3P
NP6TpH8Yew8sYTy9ALK80tBgWUt9cKNTjDZSjotQisf/i6WHD6KhFAoSmcHwOITkAMzcTHJ8Es1N
SYekjgokYyqmQOwAW7O/09ajDqZzYGsugdSd5WEt4v1qVikgnoLTMomv+wbaGou3KvlbvH8x37zC
76nxbw/3YPxegJxBdbLxXs4iUODuOdQ5Ko/Pt5Z9GPzjJLSY9AepSpFdS3NRRw5L03Xkc/VncWLC
8yx+dadqrDII1ChpIPSyOxoqMrvAnNcVSY5l8gxh/oSqkp9SrbxOBF8zoOWDsHbSacNZ10gN1qi9
dgaHYr/YmGPh4u3kmLAZSGHYROeqoBMPN4lOVodkqfFtwuSD3m1a9UwzuGVX6499Jcj1R96rCrHv
vXbTfHJQ1RUlXPgVRXEKcn2MCA50T66V3UF41EhNPx4PYwJWmxAc31PdArLUUpQONbBO6ji7X6lO
GqTpWmmLWx5QZXBxChv+53N7amSEy6pECcLmdoVBAZ4FMmcOltSimQkZV5iTg+OBVnfh+v4GS/1A
qaXQe0Wq9oJoLZsG1eqDf4aFcLThCfrXvt8IeoZl1oAx+XIKY8QUAihb0xRTU0o+4W9blbHxo6N2
Pn62CVgBmt4C8EaDcUhoEg/iA81krAonvAGRvpls8c04nKZRrdI+PzBitCqe8n14rpaDwIW98L61
Gq1eOnf9UrjE7fInjeuzG/EJmKxNbeq2I7xY6kdwNuvKoWj1l9P6o9raYvCuIg6eO6WhdMR+EKKr
NUIPmswnnfuMNEmruXXMgNz5YFTbltiTiIK1Qk1Gb0SZQYfRthvAO5UzwyHPruZxKrD4dHv/EkBe
sORuaPBLNh585qRhDdtFR+fq7e9wSh/i1MpJO20KmQDNjizjFNRFc7L7VD/+Y9Xfwx2WMD3G9fA4
aceXfkadBHJ9bhSweNxug81GRHuo3/hGNqonBNyLZagu4JHv+0K+5lbiVz2lMrz6AbwVb+JVOOR/
GWLY7xUo7CANQvMA+TMbTgkUix+3H7dG68MjaHMf4IO7l4OwM5HHrCZEBJCStFO6iOVECpFpq7pw
moGqprToL0il3ckZxcRZpb49LpeVx9ismoa3Qk8ptb+j5F0OhNMCgy4xR7tmc2g4gl4gyp/f7jE0
63NWmdpHKe/sESorlr7fjf3htNOGVXHz0febLy7VmNZBKnUqlWkuk5s4jtg4V/GsvgCtSOUCjloF
ZnUC7sMP6k91pd1IIESMK6qt+m/9FtAmphttIU7FClcOrtGFcxQlhF3ldq/g/s6m4IQY49C/dHJy
freFnoC0FLFN7tkGxepIhX2Z/myy9rd9gmWTzp5vBXn/p4o7fCwr3c5EDaHIt/7n5jggauI5kq0i
foFRQOoBvg+E6YNGKKW1b9p7ZF4Iu+hbu45k4bm5fyg0sbqdxw34SSbqS0ivVD6qWWczNLaaLUKt
M4ZI6yo8CcYAcWmF0dVs4NGpA9Y3/oFv8Dc/zKD5AVYZNaaYTY9+FuD0gPg3IQLX5Ljjx/kXXJu+
1uWAq4Cs6UVqTeCscNpXfa0hyEHkdU39TTlnBknFzBnY3ICELzTtrR/vjFgdxZGaG2V6jYT4uLVa
9sdgefpXwzRDCiTAaan3oG0pg3VeokvkevlkiIh9zAvuQi6dz7FzMmIhDgO48tWEsF8dJyjuxK/B
TWMGalnwTGdAvybbZUTFhACBcqqIcnDICqDiKpGh7gD6Y/7RbyLmz1iavCt+VGIUzC7lX/9v/Nrq
8Ixoc50Y81/KIqLNOSK5wkVezdQcfjs9kUCqR2ahe24Eosf8WDl7h+/gGk3gppLtVHLI3TKLvgNg
Px5wZm7yj+caPEdQok+zlUOlhBqO+4cs3H7ig0AAF9SSMiOuFtgALjpgzUI2QrxV8oHiyQoumgd4
yqumGXitXBeG4pCGl9ECTyj+09EY2cm/Ui17jfcuBaZHQj5dpVeNT5QBe9pfYlBZFRwh4YYRTUps
ELWTou33TxAxcd+Nc7jBKGLx1YjlHra+JcBhW67/I/TczMMGQlUkrNQev4Uc1DM5GZfKkSx+oCOt
fcFGP4ds/YLzyIwCDm5PXhraDV9xDRNgLMyHd9/d+id8Zyw7LYvo+s+oLeGHw3St9wDNl2xWfzI+
+vgEXGCj2mJcWaND8YylwrV5EEYYXGg/MPgToNUcbf28FjTH9aoHuL61mRLTCkJX/zlxGbkv7VOn
6mWJuDwQUfxmTkVZ/odqYGfIchlj37uysGtK4kg2Z2tZ76qXwoL5ux7Yey/GVmluSCpuoNf9qSia
OMaiZoMH4ZMd6B7jdNFPCVQPLZSoAMbxMSvPmQk1ppAMKTyYQksH3FnngJ7kIbZvjTIAFM3jbExg
qFJO1o0z3h1E/eCUjBOA3kvSDTc3PrwrW+g+7/dZwLzlCFHCBD7mdnVrOfL39PvjI6CLZHiLIVuf
/qg1o8IT6ihcsktEc9RMlcM534rlWk7Av+IafHOBULqENN1ldgd6qCo9nxCPOhHEP7xSlXeABoNb
gOyauMfkVdSjNI+vIhvlRnpPdDi607J7fPobevjwDS+J7DXUtmB26jKqnxpRYcvnD/8l/cpD/lmn
QcCh1LIjfPf3aZZq+h1Tlu0hMEEiq1Cf6zrGTONszffOpeKQZtgbAc22j2TWHBI6/roJpQnYqeor
RuJ6eH4EODSYclXdzjWEWPl7y/tcW5TVkp2ZTOoYtcrCn9l9v1IK5hLqm1uIqgkWsBruFs7jeCKN
zEcM+AdgCiST2l0PzBvaVwaM1E/eDlc6gLhKPMooptcod4Oy7P3fphwPqYR9ct+gGUcAmn0Rn3rt
r7O0zZDE9K9PUS4ouTDjdWQlDeXp8b+MkWL87zOQI89OpmNukRvscApk3kkKPiz/cQzsW8NatSXX
EV6qqaWLGpAVx4b5bL04d/S0vPmvu55ax9hsDGKh4cOsXl9kQ3XPBtyQf0KRlhhnSitB+hMm1uqF
s+TB1YF8wPl5hzFMQz2bctJ/+q+EUei0IrnXB4lJSsILykFra0/LEq5aUITMy3zIZGkv9z1+xQuD
Fzg+rykyqEOQCIBmQWUpfDw0uTl9DczFR6/63VmVfpwwUd08LtMn3W+asFAi3KKJQUu6hPEkXEY/
ayb1AQthHA+Z+efLg/fivQlgw/lWZFvXa0MTL/FdgsubmUKm4pcCuwyWFKsM5YKCh9HQZPX7pfLo
t6wqnrwsucgbhX+uk1kZ+mSST1Aao//13L+dUM07tArG4BfCi6B/gzUXM5WOmr8rKhbPFVedsRtJ
vMN5WMkucmK+wcK3zIjjxad203D84maeBtqWKemEqu0/9sZFl7r8lw8hBLlZOMicdiCUlA1HXATe
LndFOa8bIhVUCKG0oDNbW8QFtAUnd1/juGUBciYfYfOKOZ9qspEUX18nkArm6kpDbZ71VI+RyRxo
j8JeQIkP9WsKPclnpKOQh8y2beTExcDuo7tFeQVRBH80G7/OtZYM5mATdggs2StV1m/9P0eo5LI2
eE7KGBgUXudUEsdqczdidyQD1z4HfkRkduzQOdhdoJPc9aGMac4vn7kh4aBReFBvHnOr4gaxJQ/E
lsdBNHviRZW6/FOA3lY5e8opLyoN2vTBjRrXWdmKg5Fx+5v3+MSGgor2TlHn/OTQBYDZWvqwVSN1
QhfPsrzW0BQP0JHGOnystvN9mbFFYn4hrIxo9nPzM0FJOW9psYZjNTFSTKY79zxoDQ1XhMS/JFsf
4wHVj9Agz8aPr8NfaOoOOtwZiWr3BdJzgB1n1pfMWfPeutlfuWkVFlfiVnjVVWzYaOjiWD9nqVv0
hkVBKuDsRdymPxn7ByU+HXqD2DqR+Fb76KQ4exG1UpHsHUyAUKCHICyyDLrYgWQOX5bc19xCSLbP
qKBx5Cc5kYdC0meP03ocviOYD6ARlOXmEvWFkPBoPTdDOQ/AnTS6CgFiuCWkHcfFO4yPgLp1e3tC
UYdtH0EbE+6HfnwO45IN2Ax/RGLfbx1cQ/rNIo/ASTZkeXZMKPm36oaN0HqHY0k1wD6jhuUta2Zi
+Iow8b/ZW+A8yVBx7UiAlWwY8LnbmGtNGt4QPi9xTbS0c4ZjRAig6tnk8RJt+Zkg1/fIJDdKC3bm
WUOrCoyarYHRavRSe4cnFreXq1VQKeyP15fDwfaRnqhF8qEnFArwubH8XmTWH7V3vDzYrnd9Xqi5
/nFBiw8WIT1KSZVR4LKxA969AUi1/v/oVU1sPmqBa8qBAhh6AGkJTf56mZ3DP73kqIZDsmp3Slr6
Fzp2XpVqfirtIZCtx4UvA+k5wS2qGjHjuhwgUibcAIS9kchcSoyejtKUaXH/WyRqQBzNJ9GBi+zk
oNTG8FvzaBCaJtAMACrXmEyZLsDFsEHUYzclSi/clhtMRlo6gq7lFS/HwLt+YKFwG6m4bpcK8YH7
kq/p6Eh1KCRREcSrR94u9Hgas0JYF8uP8y8miDD7apiNo7T281GTNH9RDbmNzueNErB4LmLZ+PnK
UO73UJ5sWzOO306cFSN6eCACp+jl3w+qTgB++y3WGif2HSZBgQGppBYqaIK24Z13naObtCgJrMDk
silXRh5uTbpnM0tVLeae9M5YCVPXu6KemUlZARZajCly3cTijEX8ThP5ih/OTZVFJpeIoQsJEJYG
S2wRc6x/dL/K8v0VUsgS9EcTX/BbaiU9FoMWU0Ko1xY3Y7jz/avJRs1Q2mL2s3xzQ5QYgjHTmYNf
wr0DcArvHWIf46sk0VLTH9huja0wewH26iGBR4+Ox8DSbV1B58q2lh2e38AcGZAh1PIUh2becFbJ
aovyWosW9Bw4Bb0izxQ61Gipde1LcpDbZ3vxdZE7IDJDmcHJoBfshzr4JF8dGkk/nLqJSTNBjgym
a68XFtZ3gnDBHNTCdKkE3Zc42oovkni3nK61MpcaJC9LqfE/7zFWbvdnhLyywm8stmR2WMzilxWl
S5Z7pCW0eE7yNx+X1NKS/FYPgw5t+0CONh4r6TMtOx56kJ59yu0p1p7xnzoEPQ4tNViMT7dumShs
1gV8y+hqAG9ukUtkv2NskIedtiBkJ4MZmgvHg2sOSTiYs2Kz9Tc206vqENGBLWbc5bsoniV89zAG
IQGFF9sz+nPakVzHaXtyMXP0VgtTobmmApDm1E7arVU9FLATLRnpnxCPWeV3SIrmZDR5TI3am07o
2FXRhJUsSMoejduPjrobgsEMYhx81Jf2kOzGOtioPyX3/ZqGIYPXT0C4mltzhHxfoC5Tt36gkAUY
x4V+H5e9DX4ByJuaWm1VyB3fsBHdZJ8r/omPTWdTMcmed+azg4NZWkdzC7Qhw1D8t4Dzky2k1bGy
R3hhds0DSyCg6lYOuAU2d4UhHS3Ulq7G4L+2rw3zbWgxb8QJlLVF4gjx6Tyc9rYYdYuHWV8bLhEL
58FqZc6phJDYUtURkVaaC9p7/0v9pq7FqVKLDVPZXUepnHg/vIe8OOWKgLUlbHVcnrm9BJkBAnPO
U0TaEyEDj9G3tkpFfno1Q5u80z3NMd9IcgxB2xo3+rMmW0JOsaKpBENd8KLsVP03ThIKzOs/rWyt
C+EH86Jii38O9E4B42VJCODwM3FpnExHkIuwU+eRm8dn0ial792axx/3cXn8U9mmTVReLjm1thVl
mnOMACwgGba1/8mzSTxJn1BMbuwLOxWTX7A6cRPDIyM89JMGO0iblIfWW6Zc94ZI0LD1kGgy1Qnq
wKv5yv6rTS2y0VNj94fFEpd+7ZTtkzXYZ2H2X55U1deZpFR/UZFqfaA3uSWGod9BK9fC8XwyUDSI
BF71a0buu+k3y4PLw1EeDGuUs6S+3CQBppRrE46YyM3vAK9XpS1CgrQUdXKC6DEQdbCx8ZHGscSV
6JWu7U9K5J4F6wRprXIcKjboZeOtoy5GaLDX2fGI8okG1hg0anx/BvIPf06/tNJAX4eruiSK1T2f
ysjw2ExlFpOENx9X+iIvzt4VyM7SLW2/tke02bMNw1gMLT3ppCP6eoqm1/QOMRfQhBOGGb3iB0Mj
BUJymcqp+mX6xfUmetHIyHRMy56tFaEiWTyD7RaZ67QR/U1ylHkjw2UX1TvnBijE4NQBK3T1OgqQ
TMPyJHMOxEIsSC/fKs3bw125HuGkW/OM3eoytFtsx92EvQJhMWJ/5BKGCzRl7WDya2yJ+gg7mbPV
K5h6iqBBdonnUiLVhNkjhM00DBnlunOA+Tvtxbv3/B3F6ftkiKueKbItXqio6XxA/x7rEMs69fzJ
F3fpffoYWjMajzwNbGuzzgsyHop0ktHl/NbtIYBDSEPTXUMto9E88AQwiZfA5wdsdGWaXIYeT3j+
pek7o9e1/0CJMTE+eDIanAZoQOoqJumDeERf4a+J1IVxgrfRCQQg5OOe74p5/sDffOyFQaxPq9az
7NO5MepQCVgjUAFkBRLLaRhDQQwdszL4Gyx6GNjPmrL2tQIS7a0xYtme5sg77KG28ns2qB6Xtpa5
uDcUi4aXxVAHtQT9YpizBYbi9LCWplf6n778qcH3PV/l/aJ+lfWQK8au36UfduLA9ZGycFzJOjsP
yvvK24GPdi9KOTMmw+eb8Ba+FFwt+ve7URXIZRjSYVzcBkZBQil0f3+TnVw7uo1/dEChBWZUhezX
Fl55b3JDyFq3J7PUF50pQ6trmb64ZdsGq1SKPwXP16uSY684L44fSULfqRmx7xE1pRDFMIKuMiLV
qRVONyTEsiemPWHuYKVAnM+zEomyp54M4zaUvj+Od+UZfdsY7iTgWe8zrXW9teY0tDVM8c+X8/SX
xw5eRmspN8FzCub39xGxglj4stVfa1WfK15qDndbPCncNRxDbJi53ieoD7i9F3nOuisbJurgtQnT
qoQ099/VAG2Vl7iM/1AMvgKlOoHGq3p7LO3kAAJGueyIIH3ofcQJ28KJHRMY187JTIX+26ByUiEa
tOrGxenI14qL+muXQuKW38Fqzaao9AszzyheTSl+Ks07dDhlHH4FzwPZAPPGUefZ3tQ88rMPsf/z
F6zGtyKaUnb4dW2qeY4mJMey970cHWlifYZtCwy4TSycnKPDgnJfKWzVQRubFOfE5eXSPWQppU20
KqJpSZJKdtIYajPMaf9kIO8iLMdPSPwM+dTbpoEArwmpOkP4VKn79paW57LOASN/m9xBeA9vusxh
o71PXJLxBoVuoDFuR0fPqNtQrNcydW9Xu3klaxxZfrQtzEQRER7+3IEWv4KVvCP8MuwyB9x9c4Ml
c0bfuEe+32gtPIpv+WYHNEnXu5t4FRGmM5wdZcv89sopC0y3NocjyB5aoVqTVIzKRuUQup6b0xoO
TU6FPCmmnOpbDGuhsoeG/sF4nueSPbpayjp9VltKOoRPahEu+/GUNpl5itpZ+DYduYg5gDzFF3rJ
wyO8YX0X4vdmufOh51efZn7aojeOMR/QlD6ieWskAHZA3+Rav31EhWosqv+kjUqhYeKn6Kp2oVz1
TxP7WbtQpXoTv76OKO4mutAjfxUoqcEQKHcpLoFwhEnXDKK7pw+pr2jcoAy5+A8RcjKojrQwUW+M
NWGylT+MNTwnTR6u1gUzWy7YNfMeNv1LP18tfmcl/DpNOJ+G2IFGOpchQfU/fta3nTbXsph+Gkvz
JU5BF7jLAyWm459aph3MExOL7tW+TWwW8dlHLkEO4Hu5UrBZ7iNd9BFULK8fNy56pw4kqbZZsQYA
nRcKfUFCRpf3NvIAfanSEjXXGSsWdmLmHn+shApQ1K9hZGDW5OzZ7nRYOkh9UxeRgZDcdWXdesw8
sXeZ1/8YhErQJ/QEWlFM2dcFox1uXjbcHX6tNnnP3oYH62gYrY2UM8jubTdYFndiRKroF0HDWRkb
n4A7gS37gOOA365RLf3nFR4+N+mNdisyOO/4ShQT5YlrJmQzktB3Z9QfTSiQIWI0n4R5K3OUhwZ/
wad5iajjNXcdk0WhYOcR1bLDglsNBls76rL+8wEwmPXLr4i9XuNvVhJ2+t/xqeo6NMvi1QGsT+3v
4Z0wtPw7vOw3psA48gbYfkYVfstY57W2H7IAjFlZiUBzv1y1UslOf2wJe9GHlb1ClXIQIkCS/50/
MmofuqARdhcaovcxOwJVNm85OkXCzGQu+jXTJPtTWtlIG1X8xsxdPY7zl0Gt3/vgeo5L1rqp5zbX
DAEsbFqyfTg34HaLNAL6YSQpPMe6SBQcdxKhp+7VsdaArOn7MlVA6GBSsTrOVRaGbYdqgu6xfvPq
M6ZqSYF+qB5FmEECiO3Dpss/2bR0Aa2vO/P8knwgyny6t5f9UyJLd+ojNzVZjm1TdoIJpG7jZ/vh
w168UVc4HEsBMepPLJUSW/p+et3SAL1mVWnTUEh6VCLuOlRM2WrnEyNlU47HmGKT2ikMPU8fF9fe
UbavQt9MSMGN721HCGHoKifLGPPb1BXrvxgMC3dl1b2v8WAE8zYLnCXTYRLBye25XYMEHLZBNhdL
w83ksjWEEnMhDZM11iUuGTm5W4KSxYR3icwMJyDFI4hLVClvRLkste6ouONoEUg9y+emogO2U3yw
PZVfilUUMHMOHhUwBjl3JGsV5rU0kc5KyhkeYPg9uYSwAKxLM4ejuxNgFKH0p/egG39vPRN6qiyr
6j9fT8kvI7jGs8sN11eL+gfn5B4/GZqbvkmKSl9m29R8phWBqdqSZO36BiEnCjZz85tZ4ZjyI+TA
WwNAnCYiai9bbaPw7YVYaYlaD8J+WhQd5RH5dN9TflOlJ8S5r103jofLBGzhMuOCBuCKN05AAPsQ
feRqVh4lJ/K0lDLNPUnVc25GO8YcbqqBJMxtv7ByZZxWjBMy0JGp9xSBKSq9NQTCgGzQNqGImyFD
8f455JhkxSvmJtL/7HFOEVpMFuBtrnxmHcSDrlJ2pxtAkZFUppxCBPHhpPy2JVeoKNLGBapgsbvf
DQ5LA8SewVQx5e8Mb65RSZWYD2N0Bvnw4MptcDbEfh9M/bdA7enxbjz/e8O9Y1GYKMwb8fDJJZHv
ZVUUhpkmdFjbTGwnX8HClkssp5Q0CYLxCgpgRYf0lgf5pKU2GusptiwDBrer2RmJ7OPHyZbbzknX
7r8JHNhLWbafwOlTkvrgrKnPg3cQbQLn07fPyu4ON/eMyv1PNgmvMwZIkYVQSnqcXcpHigif9Uoz
s0mMexJZQnlrZWO18tA9f5sH7jIHgv2l/Yxo9BKtWRdU9ZpvGTaGOTe4eQmaRDmu5TobqbgBZvW8
C60lKHu4l1NHCSLq06mLXCdgwP/K1d4sEHCXn3RakL00riLGhZB6sxxWyFs89a1zQ0uNpEShyXH3
X5+PVs8kZ6tesE6sKUsiV3zj2iNAsva/blmx3FH6RSgtAiSULUG1ZSqcQ70w4b1+pQle3MW6dYgE
X29P37Qm+J7Er/8ykwZAqX2k7v/wCTGDGlciZ5WOz18pmuXMYCv+wfDgyXKzdAX+VeGLTO9nQW6c
0wmCDDpdchPsWdGrkHiFn73zaLzEC55woNSiwR0VdvalgIfByW98CxUbsFxfPphSXmgXpyIZijNi
T+tKYgasWZkmYAg1Cti8bUaTWy4/EJwWR9X/G/2SatieVwvXpagwO5G7jFSsrWS0F0WMb8o8rPBk
ej6AdPYavOL5jksklTLrIwTScCYeJyHhDjtNHpEeQy54ktVvSYQDKhBZCOhuURfDXNt2F5Qb9HAp
Y2AkpDeH7XbhCpSqQ6bkHunStF2kdXjdTHZYo3eO02Xpn4szO1k/uWvxJbaxyjrzK69sBB2NGfLj
IPPLJ95tz5RFuN1xrqpkR0BY4KMr+1hdTQ6U4ik4QWpnr5gH8ROXX/PcWY1k6l10bDI8TNAZZ+pP
PipTZa4sbeBrE7xnYkr4Dv2fbPW0Mthbd21FKf2bhM0b6B45/8JfKO4jeOBX+tuwgWIW4kPg09dT
O6xhwA2r0otNEh/QiUnrERHDxgEdnPfDsaOAczpqd2opv0sd+E0mRI/mxcPvzXRxy+459enCvdTn
Vw+JqM5R5USIckn8DgOCDMvvoSaVPTIe/G4rBX7mNXBWdD/3raIz7a3tsr4rhlxt+kKkzJR/BH/l
dN3ciVbShE6rlfm8i1r9HW7R97LcnYKFTdXe+U7glSRCUkNlvLkyexntj79oTzpWrzdWR5g6YAii
KuNLIdltW8dcAlPPuhQUDe10khSJqVozm9onZixhxMceZWHiJ07TzgzJ31YSi0F2PU+W9dYFfPLL
u1Jn8irdOPp1B8s3NHQULyTdQ+tfOKSJsQzirfDkVf6hmpOmrvt1SZp6MmNAzxV81oSCrYguYwjr
0qNZE2jo4LdV+XRSftt9p1nrLfdfMzev1EV4i09OSTTrodasLgk3J8bWsU++OlvlOfQ9WTQitoXt
QDP0Z2wF7EGAojwjl1iLc1B2FO3JRgSkobciNIrmjZDvYD8HYCOQCcMHGKFltCmvKSzTzskT0zai
qUe+emhed2XC4Q3jqpOCrecUus4/OgW27jmZk77nyHoaAuekR/dVdOp0GJWzNu1ef9GfnTgNKHvA
UGyE8hOFPQjb3oA+EzCIemzFUfJSSJ9z/iGp4edpkHtoC8lwgmVx50id5EiGwNNWTL1bnGDdjxMC
hUrPPMJvzF7yoD9ewJy8Ozgm+jPTO8dVLG51VQmdI6og5apgh1eRvGb8PmJawDG+aM9trzJtkaXD
UnIcM7s0PDbhokguZzbfx0dtdoEZXLcNa9RLfOliKsUYZE1V4JhYPguw95/BDXHfSCdi1Oem1avo
fGHsLBIlbZoY6S+amMPLYydJEJ/ZAO/TT9kJhXJKB5ZxxBlQIp3i87z23fNPni6ApjOOzkIFxrHi
Sw1KWCIdEWzezZrVFYh+9i9iZ8ixnxpA8lzVIW8q7avYUCAhzSIp9fHvjzVbMvisukKI/aTMIR3T
HObOXSzSeSnrkyhWQ5n1tsxi4jLiXhEE1Fd3RzRuD6eK/3Mu6IW9SXw/AsyYwYdtk3cyHaAp0s3r
5GEafysR5Y4+vkxUDw8YHS0z5sGqIHPgGCydZT+sE9oVvpQ4sXPhXQGDY/Lnn4VuSJpGXvJY6QqB
uEDYP8bkVsDP2xZmJK+S737L1Fu1QcgzGbAE7FzE9iV9fcQVM7D7U2l5R2eN7U+t4vsK8LW06NaF
17Tbt3JvVm+W3m1x3QnkKXz7UHhSCpsVqwVzpnoI7Ny4oYTvtJgtPOyAWznJnxQryynxO1ikevvy
ggPRWmp/+UOagw+h8diIoiApIVKVy0CivyoPguvbIDyIDbO8ZJCa/0/5BREbSczu6YvKMstpw6eq
olP5sbtDkEcrlQ8ynB2i/O3uKMtlPJCr8C59o32zwiX3Dd4Bzshs9AIWMPC7waa+WDvuiFfkpOnN
XrBzp/77pyJ61vhR0h4L0kDf/R3rWTB96eh2JcXNHPPiXbz11o2kvzvBauRQ6H2OpE69BKRbcf2t
1cCB4rsOHsFaM7TUffgIIObYaKnS575qYIVjMJKj6A4Te3RZ+ZYr5IyjB0jWZZkISZGdWYZrTaF/
Q2aRxbFV902ixSouAOF/u0leJJSsXaQqvo05J6xa9AtuaInc6F72x7COPpXNoooKkHK3ORbMga/r
Ttya0SPM0Xmk4lZNIIkuKZIKdpTZcItDRoYdaQH+P9y6A3OG8bPUQpDj4D9okAKK2K4rYpMEsUOC
AaC+VZsU8P1fI/3AXa0v4PZTkCWKksjvW1KYzzHxT/gwC/7OjIg9UkcvyrqpSero4MtV7gBDl5E4
ZClacsWfGBXUVyJ7XSZA85iVs+PXVlDlGoL1TB4uEt6flbk9awPIhKz3fRxgl05LzO+CpTjUikgU
6R9RXeI0Q2eh/W4uFYv+tRaF+IS9XifzC3imeje0FgAg//h4ar4Wo09RQBse3kJTQ22QSsMRpk0x
Jr2J2SF3rcCpNeNr6XjTDX8UDbeEoAnrY86pUQqXz+FrV96+1tnAveSaazMEfe3U39pnnUHodLYd
Sf9REGgR6f+fFUIO6vrq2h/PpKWvPQPdapY0C/mV5Av8Dc4AGDdQJWyfVQkP9Yh+/qtEqmCCvvVw
PwhWQsR0pNKOdh9nk8Q6srzgkFywj5YtrXGwwLHu64Pd0Tk6K3lYQ9MZXvLa7dtE5yBSSaEB5PKI
dTkzLMFUZXblyruby0JvBKnLRGsoBjTnGJCNZDfaFjShsSB8CPtv7WFQmrSEDTxqUl3RDLaE7LUR
vlJ2U2GabbDlavimLeecGeTTyMGPfvZRu8DP2WOzf61ujiE+FgbDq6HfumhS88Wt11q1vBeV7vA8
Cq9VXgXDi7ZaxqRERKNAlpX7/y+VTJMXhGwfiszGatwAybRpsqppdZ9EuHVCjUUmTNEJWKefIWGM
V12yqCeEfp3bDBz9yOW3lkPFv0E9qO3x7SLjKA4V4k+1shFkz5Mu3YhQuFLiqfT+3Yy5LoMLQfs8
fm6go6ph7Qk+WBofPIWObNIZTd1DA4jxqYYO/k0Yy5A7Zp15KNW6BGF7NTrO3ZWS9cWs+ySploGh
S3rb8K61vNM/UR/cs5Te6x2ne5l/kkfudO3P/AQoECjB2JSPNksi8aWhmIztAtybd1Rvcacc3Mkt
7qrJ8liKpQ3LSZkf3vgose1FL95m7zredoprXqFaS2RgdTV+bqbAQVimtf4qr5RZwyQ4G5+0Jeh6
r/lNzuglrhCuXsHzW+yIxzt6GLps/XZ+afExNucBIk6K4GnxE49f0/JhJGlr7+pMBDQW0gY82TEC
3Ym4RwkJh2GWiFgmp5HSf34bDj1LKRwSbYdrtxVClFLYIV0a81+hCq8XY/F+tpm0yVoMnZAXpCrs
nvPD3nfv5ASORdx8E8SPwa6AfbHjGgdwHvgR0rSR75kxl/1BU76hPcVt92uePzL+hnP9iCHeVdnz
F1cH5Tv4ZiPTgAiOFSouuazjRoxZm5eIff9JiOSynWI+EB+gnmScc2ulQMTGm0GSM3Z1e+0YvlEm
KiZExAFKedQlnX29iLmB2VQ8srCbeRl/ciJAdPidZAe7s/wcZNYW8U8tJ6JIT3qXVhE8lqgsqkAo
s4/osfisX8RLoYPgK/CzcpcFQxDlFBl14tuWXLazcg1LL7XxyTn0xaActozMuBFIhPp9eG4kfNld
R6KMAOlgBnEQVa0aPiwqM31Qk2s759JlHbdopw73fRiPps/ZierukA+VpCzghJUclrhxXyHZe+K/
7KB9EO+8GGIWWAZW64r7OV3rOqiN4UU0XhPNgLrJcJFboQTH/GMN0AErEjbHIR1AZmghc4zF7D9f
GRk8wtpNu8k2Ga4STyhrfS6kCZFOwAgvdCB6WACUnB0858+hLrUKLgLIyA2HQMRRBsS/xLLH+bw0
AKzuHfaLdakzRRgdbPVkWHmjNWT5VJu+mVfOS0l4YHNREvOyTWF93Q5ftM1FnNgarZ48oP4s9pKZ
0A6NOazU12OyOg1ncSC3sVuOw3qlZErKsZfRBBNdfNUgoSNh6Zts7Aaw/XGqB4PSvaguA4SNvYEe
TUCMDDhpyhlfsrC043xOWVFXYxO43juUhutrAU5fZn1Ttc1dM3BQkcgNO+6OG5lxIhJ4q6uqiId+
8l6Pv439i6G0K9S9Dko06orxUwevfr7TpzLphMEXE0B16F9wgk+VYHZoaXwFrTrDPT8h//iQ2UL4
5npER1LcGi1ebKbbv4H5QSb4LCA/xsQLN43A2evGHb7Cqk6X9oSSQzX7x5HA9aK07rRQOm/8PnVe
Qh48RacgsIxIf84KU1NjhSNFZ9j4OJGU3BcPfrIQopMDpF4CcPWDofM7b/Vmi/oCgzKs3yxhjkb9
1u4vt3KMZ7XQnD4xHFVFnTUGqYqrxp3aUQ0bCw8SYn+zURuA9W1t+61t8CctzSjQ3SVqvFzfO4G4
bJ4wBqApdkJZ4wWLpeWyrbQG6hSj40GSKY1MntfqUDhOw2hlrU1EYQq4tMrSvAO01RQktxFSfeV6
4sENleXROQ2ytyv6G7kLj3w7WfN2F+IH+MuJRsaGtnaSCf7S7bpPeMMKcw2uc4UhkN6do2tjQpMn
RQGf2OpidsieE8tZqRb2aamFTELZZdfQQ98x0RZrSgRzaBwR9wAtDA6YuVX4uKEDJI+G3y5I6reC
GA8iunh33NjiwhSl/Z43Vwrf8TjxuPSP3RMly2ESzsy2zp6SY6V52yRbHGHO1WqAvndpChgEM4vS
luMoD7A0n9JzlKl/kyxj02cl5dhfuay4CMcHmHmDdWhbcpHr0IxGM93x3MdnK2D+6PjWOXSRuu8P
GWDSLvD42ms6QmW2eJtaW1djac5rDN2oWZRHjMac7GwHrBdcASMVOBPO5fu0oRXDRNZtIQ219tbO
Sh6PBBeyxxZNaYyubZrRnTIGT5KHtiv2VKQig0zzu53u9zKTRaTYl02D0dr2P4kkIiX3AomAZKpG
c2gSNiKdOTeHEPVJgHsWLYRAhtCN+/gx8g7T4eZOlaKXeFi5D5wBnPHT/3Wdtv5w0eGersXKAnMu
JHZ316p6QNVXAQ9Va4/EmyhsJUGo9gOMmgzwDjVnjHaXT9dP6V6sJzasmzKY3gFn6fUuNcZA91T6
oUyFYFWSu91cVrzUrDhlFCYarZj7vokPJ7o37G0YvmljOcdDlk7O9bhCMdUTvqsAe8SsxyZTm2Ws
1hZPDhFzFT0qss0GXukBhcLtsrekLU/hzXYqOTE+bdE9eQop479uXNUJE+KQBNQleR3x6CTkkENy
C1mJC7LoPjlNLTIzmBuKoUqAu6UkFe4us9+Y/LhS7GzJNTR6Jo3aIxbhyYMTV6nV0XioE2cgdsHN
TRBjwnW8KD0gMYZX+aTd8S4TPsP2vFAMiQvUjiVYVc++heEiL0w6H8HYxtwC0e8SkvP4JAUQHbEa
9jKOtnpHyH9PVBcCJ7DAREH7hIRpFVOTz748YuewSGak5Okb/9HGLVEjojgkR2vtWVwlJc9ZOoGP
EeW9guFl8KiY6WAE467ToaI4IwZVdRRpElWaEElV5sFZofu3T4pkt9flWREi2sMGafGD8VeJD4e4
CVav5sl6P93PH7gJpvbU1Xebo3mJRPqo9AgkbUZIADJ2LEgCLErykkwwzG1PQEUnpHS7OOioTcjE
PBMhsTc6r+B8ghQQEt8R9jnlaU2B88wxq2Frcba0NihN3Wsc9SmOlRnrQjtZw/hj/oGGd5sT3m7G
MWHInVd5VQ0RkQ4wCiICion1SquUzLihKUU7b1Goi/jBpTJ4zqH8oo0jbSdqXcQKwQGPWTqf4JYf
duH17G/XEOKxyo8TdNmOWrL+3mIJ0lUuqkTzFkbSptGLkPMEpl13bEPhB1ao8NgDSzQDn2Gkq3jy
bT30z4sDDsbIK4qc2WZFS2czsGj2w6gqpGR7+baWmPrVo0r4tSDKSD46ozjf2+oUOj9vADcBkR5s
ECt9oKOO6gM/AeEDGhSt2rEz4+b8Uipe6l9kk1n7Vv06dFRfmkE1VXhgPDoHWlQZp2v40Rb5syLc
TbJOwS3p2IolzyVqoQrBVNKNf/NpqxAiLMeE1duL/LdHnfz8TDvxRZ8hkeyQ3xKTFToA+doIU6x9
fRp86XO3t0puN7PUq7S9akmvfbD6Vx9bMNOrKsCjDhlzkUpK29vVbLL35HFeTbpkc9vg8R+xYJqO
2egle+AuawC7QO0qPvyCT3NXxprIlFvItzgv/uhKFDTlvzK6HRZuGq3ZOvbAZ9a723fDEpa/iRvS
Nu4u9aIplCkX8EjG+3nvJ+ih9Bqqw+IsWweHSnBVT1A0ZLdQvfLF27XnoFQI+Z97+YvsSeZhbIE9
MbyT1G+lZ3bgqfDCGVpAz6KfQWGwQjoyB0XZTIrSNSg+KimK1pYQqvFhfM4Ld6fHgQd9N1YpBkA7
yrChUqviUdClL4gxtT9ZR8nl9nC/Of35Epc9pDjsgopIHyCG1UXRcwQtLQ7zQqtdS96Ab60Pycv2
elseextDynHoqiFsxb0vREotPI+5EDm+QmX0viaAHdmvnztwAl7APvukcO6QYpor9gm65lkhS3nP
I6A10SHetjfXnFgL8AQ92W1N5qpOmGmRAQWXnRLlosGSF+3LVtk2ot33WEa1b9mGVxrRzjHUVTcn
nCpT79Fz/OazcGB5TTSYM+q2nLyXab5Q/4RXj5LZXWtZlniSU+5jidb3stqHiO0c1Q3rF6A4mPSf
O9PRyU/Rmn3nWJWboZmw5e7y63h+g6NuTV+KmnIdqQ9trJQy2pFhcuid6tEWo09WltiLb9ktt5jp
W47f3VpJpmPEvM4VoL+N7P+r6DsP5V6FpwuyspQkFMGLUg8RppHLFfeaCbyQ0wMQKvkitP9Wbv8o
fIeaeypbDO9IBpui0yywzl6AfwiK+J9m0h1NljF1YEzg1EIswx/NA18iYlVI8/5vnlCHjlbnyNre
+nbFIB0oId1kJuVR+qIpr15nUqDjhmtiEV4OeWBqMEk3pp7sT+Q/gn185h473K1MgQSbDYnMtMtx
Q31G1TqUxuTSqfnM0X7n7cXx3P4EtobGlOe9414n2CdnQCZ8YU8RQDN6jhcO4pvpVl4m1DNrZQT3
OPiWfjKKoQUFP3AGzzsR2ccp+ZKmY3+GGvkI5bMJXr4MluIf+F/YAcua4zkkrADJXi8WkWJPV2l3
mUr5JNqZb+TSjE1jQq7dW1L9tgoxemJYwfaYtSK4zKQVinRCElS34k5AvgWr764pgJ2OBsrtNXaO
oLa9LEVywB5srtGV58gzuJ8s7ROSydeyJb5sLUN3YS8yLJPaOXvLTSyjxsLniVDAYHzpLMYpjVad
YKZFwsZZv17NQXzpt8NKy2byuaQqoYAAkJAwWPtWcyL+z/TunFPIDllLe46L1NkZDKbZ83GxWLHm
bHs3My1IUOc5T/2yRGsgepY38iCuajf4y86sYDGZhMX77U1l5zgvASol0z70x7pkUlo35w/sajWo
V63UBKgXLikEZAFs82ufSvU97GcIB9p/QkM8AJkosBO5gvVwOJl8BZm2SsSWiU/Q0ERXNaePEO1W
SclVy24FX109LNfDDi9Urqn6aIlYY3sCqUcM6tQ/2dy+1sQshVXVJC3LI/hPlOpmpc4V37n4HTcE
SInfCWe+QA5M8my55LD3rDxV0jnWFfFxFlXVZcUp7S30CXui+7+LGBTqp2ZfcZtGLc52Y/XiNFom
y/z/67QCSNXcvy+8eULbv5RCZt9n5Bn54909zeQQLkhrqI4BoPfxFEgO0N2sQHvg39YJx6GOxtIi
LPUBV/+3b6cThmjtPS4aHvD9c8dFhqLfywiSFOEcpg9v2M9/3YUYwf6P2jEV/8Va7PL7EHVLjaRM
TB/sYwuUCtmIRTAXZlFZh+X+mmLuYuTNFuJMmcYTffLc0ayOs2j7YNEnlnL4yduJ78h9Qvyu8/9b
fqoGwLQwg8A9TAvlOqs8tCGe1YEU5Md3UXwqaiJByBtBbaczSLyKL2UwQkoSpBLcwjwN6KjTQ9yf
V5H+GIOlvI+xkewFB3JObh2zJ6mJnoDzRjO/+8ku717ZT9/AbLX+RY4QWwQifIWivWGJseEAqsFJ
4Muy9jjXXo30lJAIjG+CEy1jKvM6zKJOPj9banjqW+gv38Flt0GCU6Kwnx3kCTVrs5vzIIEaKRZQ
ZOEaMNfW8At5vQI9UDAxSB3pKdVMx3oBZQ0A8ZtP1vimHnJw0kyA1VN+fywE8gZoqjLooui+IEOI
yXU1yZ6HnVUC5XWlF62jMtKSzPK1A1huu/OdrRu7bKULHKkgRuQrmv+vCd/aOPsHJfjikcGRbEXi
A1//RW8X/7LVItkdnNat7iDYLcpmQCLeAMQocY/WyCCvglxXb6L8jZClDtU7i6mdGfEhpaCnSjq2
bllVB7AND/FdRdBczX77AL9Q5rueYKw3zskAXTxsupdwOQsbB6Pg1M02wRVdPEpvI0/AvDPHdQ4h
T8kql+d2SzsKDxXLkN2N0NHbJyJAWrn7I6Ofcs3LovD5i0Ii8WIAtYJyOXrl1v/pQDpdAR4wq7rW
Gmy1fp7PNElmukDamfpVChKG9lEhujgR6NE2ngu/TTgyuBEGUvMCh5AAh57SOuX4X7C+noNH4ide
cKQw4HbPfDthEz9bkBShcU1nVcFbWzTFEfQv1kOIctAQDT2GKb+kpSLUReacqT1QfZ6zud5jAZ0E
nDBS9D5ojaiCu9pHTG9xXBJs/f7+bAYPyYO4QaBXJVRkzlCR2NZNO/LL4Ed1VNLlhspA1E3ivVsn
ldcMep59CnA38d8wAz97HCiWPoZ7iGQYh5IqD1y+NE4pLfLkYHfMe84UzAhDTfL3lwrJhq/0C0CF
HoOaTYxlcBbzv+Yj7gxQvH2DGXLUHL1H3516uF0PNMPquKDNSfQGtIA36j3csv7FQ/6sEx3XI9b3
cwCJ1MyZ+0Z8HPVujUjVQKA9U3bbdeHcCneMijpWdrDeNBFWTh/w8VXq5FWGaYPv048o7PEHJpIn
20HZ8SWsNo3mPZaBHgi/YjUTGCRxTnBnc1gbN0OsbgvpQcPkn2ebuJ0HMIIiRwkp/KRzC28vU0cf
GSTY67WeSWn/yAs4OPwOHhBgqdzPOXpevSDONaGHz2ca/2D0GmZuLFQsDAHzRG3W8rnHTYRrhYCq
HYQxW1IKkzXqU2HeCdGzcSdZNiJFxf8RjScLAYq7RQNBXGCk44bf1rO39RkouOoObTIS0d+0KZKp
INIvJ6z59B5E2DVYNdruoLfvNOJouy9y1GBcdQQb9Ugt80Csb9TEhxnQjx/dBkTp7Tkb6ig/taBt
df/VKDRdcj2F9I+jvlopwht3KWXXzE1prSgIk7IgzC+4qh0toZL8FgBkO0woKjlXuBBT8sMY2AxD
c0NXIRGMxqVZfIYj6dD+VzUyiSA7+Qk+VBg9K+VZzI2qS2xf/AZf+V/5i7l8jta+Rzhj0jXI3xQS
PkKSAsTmxdwqx7hdO6jm39PgcBOiiH9GwQpvVY5lqoJ0cMEdOMZoNUCp+1/MKaoMvbAb76MM9emJ
VwAihrF+RuajQUXgOVpcTomWL18BYWqPPT7vk7C84vDm9xsOAA+0sDl9a1EzVmDCqftePV4f3ZP6
+gs82YiTqcE6lN/uFFOnYDthqHSPMO+gdwyndYedVZfh8Qee9Q6gvLf5KuESl2OFxJuoj9IwmP4X
PS3ccEH1gzuqsns8K4Zk1OqkY4hk+4fgGbCZ6zptfxJzf80T9qdkW96SxcceWJbXVxZ0az2T4nZH
BRKZGhXIQYkj06QR1i6xEvwReBCaWqgb81mG9DF2d8ITnjnYm/sy27bzJo+YepGKWGG5djTMjFox
4Tv7NUUktSMMBbZ/8f/xlyjVsZtdHaL2kTrXK4EarwR7GSo1xqWDkhmKx9cDJX4Ta5lHdPHupEqr
yn15p39210m6IjocP3L/OcH7LEkxgDzYUZ7rBPYvFBgwSwbrBZiLBsKmvyHUCEYjvYnK1+IzeTfv
lcNRBjZExcLrwlULH/74V+xkGfCr37k1ZPZBpe0DDYWBZF7Tuj/qDxoTt7RkRSH1DOn1j6WVglMd
kOMKLmmyzIr1UEb+J9Ob7bF5+OEH/B+4f3g+MOsfIBFmCj+74cdtTjB2tWLkycnNVLEo9IsFQvyy
8EZ0sjms7jathJ8m9FJiCidORnpk0g2JcpQ/puwz7YAq6iyLXfy+fENvMCviZ5p/rcKwnLkGxG3H
8i/QQqa9TppKkAFEU+7dWfQ7Cm2uETc/FWvi9Yv3WrFTPaLttXQHJ+kIyFqLPxW8n7OF5Ejqi0RW
m03agxbpz7ic/nca9jbSffwFogdcYfx4pQAd/ytTa68JZ1OyDa+l7nXyh41jzWzDZwZjgmi1bQ/L
8dSJvPW3TAfgm/4MS5W/o3e2d43xvz9EyK/GV0OaggDfi5ngcKGJg5ZCGWaiApve4dXRTcUmyQND
r4m7HP0U9krXXUAFXjt927YTIK/SX5NqRs+L26mvwMlU/L83kFX+I9fLOAKqJVsC9PO6boO0SXix
MsAn2uTSfPLHKTa2kyd0x86IgtkKfqItln8v5gAS1T4uaoV/9MuIOY/DSdGfbpnd0EUBMm00Oj2N
VSjBCcwvygJnQdnhMIjuSayNNRU6G/EZRVNK9u41ZQ4kIaY+qc1vhHsGFwn7wF5pR8+0E30Jowgc
57MhoPx06XmgRXSj0Yd3/Npj05FGc61AUwKgSI5YLlBvVrnL1YgmnYMjwMGKfS85b1WF9AxF0Mo5
NXupmbK9aDKfg4N2VQbhJQovFE9bsa/7IkOL14gjyO6un8gcK6gSstr4HCNiUsaUx5VqJLIX5/nd
bqoR8/QgWCQ1DxBVnUNgjlQb/n0GnZImuVadZRvtVG2JAVoXlBHUre3i5t0cEFRaLNPMhC5334+k
MMltTGiqUiatTqfTiJ2V8YKIpukW+9r+CuTdsIAqFwI/l//J1i5glwvJCk7OoLQz9VzE8pphxyjL
skyZbvXv4JLPVKYaFXTYfO5OdvhOgnb2xutmXMXdsuOhfGWeUiRhKDI1zmIOO9KOS2/mfQISKHc+
rSIe6SzUMYHQDH03lbxbZN4KwmzGkmXJE2TeRUsDyOlpWV+Q8MlXQAzXRlUiSc9YagXraG/jGq0V
qf0mLJBdT+Vk7gZb/mXWZ96IIbBTycmXeYuHDRlBuxxFs1yjH+JYI3V3vDU1AhMhvm/CnQ3qTX3W
LTHf2Lj0qqtEqBj3MnrMBbwY/lHDwoXiN3DO4efaxAww14EPy+f3n8E617DLyz59QgYLJ896bJJ9
VIVD5j0/zpkz7hbY1xWy2hWmnkELrl6d9//NF5BNqG/z1MI55PFFTsnKN5axxoL2F8ic5CeIUcEn
zrPgQX13K+nq0agxt2orDkXWnizp4GvHr735pqnmETiY8kOnY5/LJDoxdEKWRDHlbY+LYsMhNUxl
ZcW0MTm0YRjnWJFzRBxKj4wdqCETteEuCtEGj6TyGvekq6T8MYmXTfv+LGMLt7x4DfRXYqyDJtHI
2bhXClWWi1eNdtef75UIlZFIV+n44PB5okQggi5trE0kK4QOzZ/bjwFs5fkMHrhHuo4CpRB6SKDf
O6ZTaYUQB7LK4viosOAqaoGpmOv3Rd/EEN49cF520E2XpcGGnFR8843o8AWDpO4MPJxIMdIQ2D14
a3m6ORApo3vPPacEPyk7hp3kpee5LqGbU3H/KKxULDt03UWknRtggoMDU9PebP7c4W5Xp6wmgLkE
5zAytne92vEuVBz8QX+DtW6KpNOp1zsqqGcXn01uYyKtZ3gGb45fEDEvMoEafDsdoBRV87/4l8Jv
Pg65v/O3nSTitz0deVie/tPQ64D6hdTaIjfGUMFSaVSwP+XYXp0zjeBV4G7hlpPcN19uTzbgDPbB
g/0hjnaygw1G03L7Vv4jGBy0s+dl+VJyXFXCOxOczOa3mwX7cco0jia6SY+o28ZtwgzbSzh4QDYZ
l8HBYIsmBFEH7mtldw+LZR8q4vEmaOgsulgCX3/k+oCwNFDuqVR72AUkBqbPCNfY4f+c/EoHsLu8
RpiXClaA0jhPnd7LHpEsQeiwxh48HBx6d/Nn9cxYUZ+36G/HbV42e1oaA9e3cN768ACIyg6PQAHB
FM54eWZKEo6NjuL42nG94VgYGIcnvpHoWVvmE69iWWsPfLzo9/+S/Mkt0ePFFJwd/IwYR/q2+g4E
ORkA3bM94p9Yrz7lYq6S0njGNC2i8dDf3fbV6o6yztS3+wm4mbEfER04uFr1tqjwEm604gXbVukn
yqJKHFSB78Vj0CfAeRgwZWnCuHzNgDvVHGwuAm9idSkUVx7Nx9sHKjoJAoprA6iJKw1dYglrgZ+T
eJFsUMnrazuU1j+qnH+LCi11zqYeBQCqYKhc0SAM6d+XP64fMt5gsc1AgwD3X5Cc6qljfC22rd81
ImJNfZcNr9yprgcJPNuma82i+99F93TjoE4j5Q444sbuAh7UROhnAdCPHR3mq//HErnx+hkTdQS2
YbgxLIaU2YI74oz5CyOoEZb4j6D8vFZ6GZlpbcl/t6dUbIKT1CP/1ocYOF6iGBiw8W7wMQd0S2Ty
shMMK6GpxKDX+37ORVaguGCLEGRvNo2yclbTemzUvBciUmzhbDwuB9FuPgDwt0JhshaONxs7iTlK
b2YO+zPdiQxnONHiqQzTvCAUdszXTp2EFSGArpzGQwmjEGnk2u7yCfrdDPYYEvvmmBw3mUeJu9Is
1GllQCSRw67ird7WsClTFekRCN+LyAdig6wAGhUaSHWKzuRGa1sgqAXsC0fak4FcxBKOxCrW86MM
9pVhSJUyTWDN2J74gPOxB7sDvYxq11rgV/wpbryJivVbvynvZSpd1CUU/72tbBo9awPxRJlVSTzf
AaCneQ8dDclWADRcCmNYRrkEf4WS8CQPD7BNUzCImsZMYMx/nCf2lYwZMx+RMx/oiPcjucixFbdI
OxgY2kz3DcABp+TyN/fqArokYo6y9q6KyMyU70hZxF7ORWjDwzJf3ua1/IfzxGJ4gXjrwa9ym8pI
0dh2LGU9ikghej5Hx/azKrxa3lqzdVowRaC6732lL3DREKYewecmgydkl80B+H/ZJpf/Iu+oJ7R3
rbeSx9pV4O4Jm9tXEwv3WFraiWGVM8J2MiK8mDhJMUlzvGL+SLETgJteqeusjJ3x67f3EmAlu9Vu
Rh9osqcToLBV6dpG9W2Z6IwQADY1DxDFJX9lsyT3IcjA0XNzh56A0WWgMpfxsRf1let7TnU2zwB7
DSzA/dw3DI5hEOQsHcL5NxP9mZXzf6Xe2ZsshRLDHvgePzbRFszmwY9tx9E6U3cDKa82+e32/xEI
LPbDKbynI6bvtoLH/BN9HUu0I0dEAPYRv40qoMqL4wrUsahSbEFDf/YwRqt2hF4c5gEEUyx420q+
VsGuxJiiuOCYT7e/cUKiHi3SU16OMqFhYsMfr2HaQ6iW1DEkH2GHN4kitX9V1EDPCalFv7MmoEfo
A477G2KJzU5g2dQ7LmpJowHw4iPisDzGSZXw0mUOe8KIyoqgm0VzB9JmA8/HfUnKddn3xXY9ifmN
HzNYM1/iP68PGz2Zbxg4Z5YTDo6wlQhmKV4rDS415oDHzdvcobHhBVTdrT2+c9RRFjpeA/1Q6Ecu
q2Ph26OGtX/Q4vq+V6gUrVMI7HeiBCevxuT8rwF3wKR8E9ve1iyi/wDMGZCbmslo1QvdfiDFN6Uh
bKdsAV1oTiNHd9Kpm/y+kVi8ZCUKLF9p6cGhiLRAA4LPIcCfl2cDekukcjPt9NVmPUNdplB+pzDZ
e2N6C1pwW/mBZqYnxActzhljBQevo7sz01snZ4rVK5aJ7eOm5wXox/l9+uW44G8kA7SGqdlqZALk
OYs4zuh0GIE7O2B2BN7FAtxmGGFlb0v/3QqRihZmaxqsXQ2n760SlG0ohPBPeah4qOeOXwPVCSjQ
+h1cUkxj4tUNXxPX/oacjtylxUw8K4+wILLJtLUeZwEJ1Y3zmiDNyoddfhhKyMHpUEI4JEY/qGvN
vBvPxj+KhW3kkS50wiYGD10mhMzgv2Ql40ZweA9/BU1eJRTIjymVmtw3TYL7vNBlwML54xnpNqNn
EZjz5UkH9esVE77rfAyLGBX2dhJ2vTmi7AaipXorEDYq9TmuQYXOu4OUqRUM8q1IHoaL+FqrI+cT
+sCZn200b8dkAfG22MixJFzqfkm4UKRrjmUUlOZRWbSrvB9BuuAT+GE2yDJKI+02/hZ7mVhg2Dtx
3j7zPb0Og36DRwLiyabP8qG6F/sG02lLLUzDOOa4aVTS6+4efi1j8cBVa2QoAY0saTVC6Uw2kRYP
Jasxjkg2Hg5Y1dqGD4aL3haYl8I4lD/zP5l6JkkFZ4TGJP+agpKN62RWdXkvdX92/+JkTP+pjasF
lLL1ZF6r8PNK96/ycR5dNbRqfIyCoU9LxnhgL0g/dlGm9Xokyern9ctmhZ6nMb3aF15WcmoulS8A
DgGvCHYdi8bCz4ohgKNITaPVO6IEVyVT7SPFVGysSisZp9zgEOZ1qkzf+4XHnk+j68+JXCmzibRj
O3dt2E0FJ9+J3Bkh3wda9keaDZePTX7JXtEtmlmOXuYXp2xmzkq2viiK73wUlUhFRoOjboVNZluT
3kYVRa2L1GJjD7Plz+wyZh7xClCeAAUOQsaRAFumgLqqgPNB2GGzgkUiT+JPFONIMpYFLD2pNQhy
j1F0zkn6KG7aJn/0PGHzTL52iT23THyib9mF+fi/lBYpx2LdQz/fW/nMZ60UUjWiq6kY/U0Ti4GA
4nyPR+mmLJL6h5QbY6IkxOfrcVZWCDwDJvZSau/CSOreW+3h8iIxx+b1KRdEi/fEO+KpPmKDjwzj
0DbAOLj9uBcPc4shJfi/PQLe99IVgP34YfIFnDfT68Mtr90vzfP6lO0HySzPfn0UFU/wPfqy/uj+
Zg7ut53bbAF5y1gKHfH/UhIXdNGSiCCBbbpc3BMahK0mZD4jRVfPa70zgg9NQGOeAI2SmKMdOFCK
rZYY4izPDcjc3fpd+84U5J34Rh1pG3cMal1/xB7FATlWJaf6tSkuACT/WDIFTuuMkcHLgNy0pH4o
bdpURUEel0niQ3Eoju9RfzY6iEIr0vyeIHt9aFXEkR9YuMU9gUOrx0rhPss7n+v8rMgjllpqR4IM
dq3lVRCThPoXwLmsu6IvTYDstEBRN1tyRnhRkwcKA6O5DGMPImIneU6Yth/bXiGaJf5EFifwjiul
vIZ+1qsnQAKU/svh9NKvpLdVFS5GKeQk6+irMD3xhfnx2nEbeoL6lIZM1DBKiHo2N4rvcI3h+eWm
0hIJdMaiIHun73lzCHJVC8rHPmUs7X/gbOvzmNRsWvOfpKGPP0Da2gq+ylvQ1OOf5gvf3aWdGSqE
zzA1QnMFCiVAGWfjGcmP6yUzfhetmbOa+qQwbMtUGy2tX6Hhz47JyewwD6wi2oWg2PWN85y7HNDF
wY793Kk9nqQTf/nu+PC7bmuV5iGkVqAkkNsWv3a9UnlCr1NJZaZWUwdt7le4Fhx8s0qOS5ehXUdd
pwBgbdsQWAz2CuV7UMY/8Px6ixft+VXSkQYuYaUiK3YNg5WeSeGtIaP2cfR57I9E8MXYU6jdLGBQ
ORHTyBWHY9/4CgRob5wsnulb030NWFRbyIBQ9+2JR+tQ9FQHuM2WwBBdldJoTk88PSuZ78cg22Nv
1lf189D35uS6oydexXIsrNrXUHu1M85IKaggMTGGOqdUw2U1p74e2lC8thPAVTCTycEjo89Ttq7b
yUyUISjPSj18FA69Ku7MIzydjeCEp/csys4+bvpiOLnsxmNzXHV5synV+E0DfDzrO1k2jqtbWTKd
yFcrupYlj6Ywvj8XbCOM1vzlGPNKTscYW/NNpSDMGsoAdmm/rkmVl8tAcu/5yu06HY40zMOE5RVW
9y2JqmGb4ah37hfZ1HwpJ2VBxdv49wWNyO2NoSFdDsnJI+2SrlSBjSv/UIGLpPNZCX1KoBrv66dq
GxXaQZ0sib1n58dFL9Jjg39fvSNQYJTUSwiekxeb3R2VYtVTpsEErppjLncgQiG1lrT8HF88EgGc
4PoV2HsnCdty4tAxH0AvnKK114C30J7bu36ytUPWG1/kc9al56TMIX0v0TfX+RyVtl/u3uDjpeYG
BqqiQGwk+C/2TdPLMeUtANnqPeQ6gzNQ8s+pQJdCzmlY9pVxgW+ZM0FJi2/Lyy00XWxCpE/ylVBF
naE/Frmwt3OEjgazuAkppV25PL0gJq9iW4qOmISfhXG7KqtnThlxJgKRbacrJd4GkykBuKCw5PFn
tsX+AYwizkTJmylNWgFlSvcnhq8aOtBBdZ82IFQTYvD6KvWwP+qvkDC179eZ2B+MHcKTjb2YFCYo
kJtTWCO3qw4jhrDDhqBqLnwlo9BxYCudPQNPppBxSxuSxB9+uWnQt89WmIOfnH+sj7DKroJZGO/O
EgZNrGDFX1qfL9IapC6+WNlTH1BKxlHMyvyV9ezrqJ5nwA8rsfgq6i38GMONCV04DPlmucwnl5H5
tBPX8kJtDZTaAaS1hbETOkMlykZBee22WfEciTkPNibLBEgMyEm/g4+mq30KoUvTNBsWO/ljDZ1K
dgxH4B8FZgmLKt85XyBFrweySBHzaZiPz+lpR/zvo3y98yplFUliIwtPevzWJhF41qvgKYjTcy/9
SAJFK2NXEpsVLFytn3FoYBthCZtMIX4UrKnKS4OFIKJA4R4bxsZl7Uzzgnsmp26nCk5MhHTX0MF6
JJ+XkTh9tRa3qxvqqh2c8sIlHMiu/PPElaY9Ao86HkypKvk7pRx9wk0Lr5r4vT5RBAVQhf6ro2S1
HRLNojMZPgOmC9KlP2Ngo5LBimy2NXP1ZnYa8Kv/SO+XnH4bBiBA/ld8J39us+oAqZmsM8JaAGE+
bbUw8tW3QbR0H2lkrYAJuRG84OZkupj3+WY7cFlQUkU6XN67q6c+YYx+d97K57fs9nhwVKZYeVIk
nmUMgHy67kMpr1NT+677QOwJoTZS0MUiNPofSdOOxnrlZ/jKG+bXCsIQuPVVE1JfyEfDP28l4arE
npdXm++Bz49eqmehZEHOTwtR/2mkCCMi5ed2/SONCfZE+D1RVCI/QxQHIoqIIlfR4FRHb2YX50g0
wtkjHP2kKitSwVJ+l99pWYbDuFk170gg5WQw7LwGRBbR07ogLLj5Lq3cuHK7MCxfXHhgKbDH2NKE
rgjIk06RaLnXTObnWTZ9/JYP/zxfmicV/tdDTq9dH54SF4E+kZ4xTRaXPs1QlfakbDNkrxSkZGlw
TycUyBtklsx6xgsm1ATuXXR+Z68piXZsWij6zCxTrZisJ3JYhiJPTd91lAnXF3sSkKUe66k8lVHE
kXlrbr7k+tNDLV2+eOb9gRf9O+67CioJpkmcI4yW5QgqSt3g5G1rvm+RUyFKyqR5FK6WRnnyUCpL
y8eVmU9dZ0tUwXkUx+ScEI8cnn/7sYNGTt0enPqbNib0ia59KZbFMASuElxIoNk0w8KXh8DsT0Xq
+WGiw8ku7hTS97LK43f6Gqp5RYNe1Rcl2RFv1MuKICkh5fqPqAnxsXQo0RN6xh99JGULNF+fdxl2
oxsqDDMgixVSiS/x6LTOZT+KlihmPSycbx4zkGcfLo3ibyHe34Dt04FTVr7xZVdKlEMUwlgdfNS9
6TR0WI8uV9IMj4YbMU+2m3VCz6h5hdDSUUQZ/c1VHeU2Lgg2LBoyZdYHH3+7m6I+7TjIVu41jds/
LRm8TVNm7xO0MD4bAfog+M82QnbL59UFHQ7jisgoNcNfDTMpp1ZTygoHZIDZwH15+MHiSrEkel2/
KUbZ1+dHyvua1+n4C0aZlY7haxFfEavV71rjJL9sCvkKnyLmzNNarUB18PZERU73ApcF2VgI+3/3
uFRaSIp4O3kdnvKSvJ0bIvtliEq7tPGy4jtlrNk7E+Tlkm472gP0euNy3FRXirZvmJWnujCFcAYM
vffGdBYETpBDEUg1cLQyLlgqqGvpMH1DWfc0NY3bcj1+bWC4V7KtMRaxF9DkQOdAgSEgh1K1XmaH
4pzULdTta0T3mcIyDG79BzjfuWdiZ7XpgVmo8sLIGuxx1HPP7oR5UNC1nbKwtcHtT525YWrn6mym
fVd1DN6OnS3VfQKCp7auy90u/JAD1DCMYNjfLC3cErPXDRVwMmVfzeI7a9fhZwUigRTRtETo2svw
jJ8Fn0B7ZosB74nxDfY4QTya0BLP629prWPfRXxCXid4bIHM+3AY6UsVvOT0RppyTBRAzyQH8EjF
eMdOspj6Mf6hAufAjIHj/4T9INlRw+A9RGd5O/ynO2bBCWiRvhhn+qh32/meCnUbOr3HkPZyNfg9
2Ze1fPBzki52kIxPnDtGR+p1xrYrNlXKGh1lc5ddiFfVH3D2IaNH+pmU5r6Lfowcod6KCv4eX+UP
qwGTPnmoi55fSzc0HqIbaC8inJW8G3NrlMjtNiYKeZMvdi8wOJ+kV2taoVAGpvRbtgiXXwy8TphD
dWBhFVbfivbzxYt8lgOJFPJ78prwPHCLacz70dxJbxU0YoUC97wCDmS7fT7DiecRURI679VFBWOA
KpCW5CnR+X/eQHmOS6m9mJmS2+hM9gQfhDdSbnYzEW86eLrUJqqK09S4imQN+PLv+2G81W+Qy8cE
Jda3ek1gfEUO41J/IQaDpPStKcMx9XSIdWuGxGagqcI1mHqUi70DTA3nXaef3GxxpHSHJs/pEKyu
ibuzByNnPe4NtTwskJX2Y1ooI0O7Fk3JrQ/m5wD9VQp5BLPAXnhqkX6cFo48hObp8zMVBrnzoAX+
afj+aq5riTPZTexatnsPJm9FuQ3pw+J7iK1GDxetqCmbwm1fHUp0GBpO03/h6uxUSRMDM8bGS4VP
wMnq5k+8kNVUQBEas/+x3c6WN8Yl9egP/oreWYMzyHO721eqvm1nb3SjVU4sHtUlz6L59pjUqynX
NNqXuwsM4gcgCKL+cIVSMupa1rELTyVYQQO49yZNIo66WjvDrcqbrWM1BNavhHsdx3QRugKQXajR
QJVVdHkYZBMy5vkvnDjQxv1shYQRAOc5huo26Pf9Egfx5qbrrBmcdB6l9lxIrLghf1hE/iqMnqdR
BxZbvGeo+edoIlaXbvqq95sLCmAg8RH825OANRsgzXUUeo0weWHXIIyxtgsw2+msWL7sFO8cR7lQ
9l/pVphSkJftOxPfAeLoqBbgLg9ovzJ4usJnWw/16XN5MMhggOEU8/MTtdBuwlaIVASZncN4d8Po
2/MMHAVZEcXp3PW+IxO2GwAsJNeGzM4JOEKv1r77S0NPm6I6OhoRYNrHhzLncJ6yLUrTboR3Yv3b
gc0HBE7tqDheLB4NQymsuK4B9uNgRWNRsMSgX6t+ZlqXMwBgDTQYYFN5ACc53Ma4w8Tk1Iq4XUxn
mxiJTTsAtxLI3q6OICd35jBkvV9zr8bJ6CJYMrCzluy0rSz4Ug1X/SFTLXq8UVnQTGZMz+cFC5tC
bmPLU1dBf+K8AtXawnVOSASrKaLxaF/1IwJseQ+KIT5EoUPXshRFLXDEXps+E8b7/8P7ejChVg/D
iu5KkSKr7kPmwjXoqSTwbuHBOwEEEdMDZNnu2cKW1oF6AoeoS51qyqZL9VitvN+rS6oMeI/7G+uV
ARbr7ME5LAC9HMEpo4n9Kbyr1rseqS1ZhQkyNo5Lk4z/LryaDWikKbrKL04d9FOU6BWyFfYl9M1l
Hw/VE8lRSF/LN1F+gY/YbIQd2uOXp6kAxx7ZN+eo90P9LfOmeZu1h9vUYFmkO+FC3tQxpkBdgAsE
yh3cNWQ1AAdXO7/8ljv699U5qcbZt3ueFUnzN4sQK/y11mPBWTeb79v2pNRTiQ3h2U0EQcbQJ1Ge
+xaXFpDJAmQBBWZaX4Boh2beeUA/CUbebgNDyFYeNOzuARBlKi17h2Yt5Boeh0Fh+dVvPpBZg5nb
GubSdMvr0QfaAqeIyg28aVjlZzLHKIW5KRj7azgvJjc7LDYz4GOeuLuK2G7/YR7vSsXGxyouyzKJ
Lfm3y4VAP+mfCe/JkkULLcFmuyG8ABY6mxe5v1GipW2/n9Rlyvux8VHFuiLZoJp0j6+sXQVxU2LM
vL3toFEqt9mNov/ckyS4JbfQwlvo2yDRVr/tDGl4jsnbEkaRKrm+wVRO2Qj5r5VTGXAV9V4eCiAt
yaCyXDAy3BDYC0EIKc20F0W85+DosAo2PZbkkAPWSHevqrSo7wFexsqZV8kwhNwlG86gOE1KUU6W
xaaqSskA7wOXkFODqrusAhHvEdykZeLYWQw3tBf4EDo7TnC13Hwk05aZyoY1mOvUKJNOiB4a6irN
yKv0I4gN6A9DORdHeZeYcunKBFg9uNXAMD3pypsr5P1ESbAWffFuMZb1ZCnRV9gPbvgXHddEIfLT
WjP00SeTyIWXG3Q6HEM3V4zkRfaCRZhg3lnBINudEYPymvd91invCdbdJ6moJk4PbM8/oxte319d
7ba55BOZJqUIDNL94MMd0G9+XMfpLu5QhCCB7JDmEfI5oIRyutq+kfBcDK0aarkrWxsetJsWcaw7
OgQJeL/KLtJhGc2MFaKwxvEXEQdQ/g0xlwxmeIfg7VMbdzXFllzBsO3CfuaWFmYv9aHq3Qe2K2gX
NAdEafJNJOjIwkqyjMOnKc1PlFHsBrXpET1/LRvGtYUOTEx/jxwsi4X14kpdcOIHzDMBNmpaW82B
DASY5tj1JixbcjQcTFyMpCcioKlx0GFv+L9BX/p1s8A+Xe24FDi8sL8SB5WsZAF+IxF2cWRuf2Au
smBfihqcyyRlXaQsAip+NNWn43MDLqZE5qULGCscReWk0MxapYeZopE1UsYH77pvnMUIfMAjIZ+k
qGLq4Ha+AbboJkRrHth6MEP+nWSWxhhztvT7pEIVjTcOL88wK9feXFhi/7j91CRs5aig4pheXa35
6YQLT/i5OUEFNg9XPCDput2ZOVS5Nq9TQzPvDj5dx5sMNs+83XrvTlCvdKU1sHP02HO6uQAkRqN1
wiYhcdnbASMnkF3t0rDppopKJ9kAde8qNcAFuMUNlaKaOV6r8CwpRie9wZTb5SY62IlT7gNdkQX5
1+HCccRGk1g4wj+1kHnpOgnS9vURW5mQkLMa7FGZwYqfmOEIrPupoAOrdrWj0EsekqUPWzCPwDVQ
A4A2fWo8hRrchK5KmFbjQhL+RBpxZGChsJ+ueKNxbBwZqH95cjDjqrqlfk8tLh0qs2vBBRNbS9UW
AzjAk4oxwfL6cq+839KRpWBuatQdVD3wLvLKxH0TN5ey55H64pHwu8zUxNxM9ef3PMO0qw8SmIa2
me4ZoaCcz4xoWOXD6GNRXGqfXw+MAQSn2TM6QaLc6utvljxiYmLxQZQBDrn6ubFwEGpCPaxdV5+k
YwLd65igYhoJc67YnoL4fMFKHXYcjJrfRoGx4gYUpyuPzwsAOlc32XY9q/Xm0dIZEQb8kt8skbIm
WSvcqDe4mXASc5FuiJGH0EjQSAV2IK9taGfOYAvR49Zi39PVXDweBybnwD/0Y5xyoQpqhANX3imU
CX/4YBD9l4anu1qud7+ejQu/Tbc0iw1b6rnjFQ4PUwFqLWWFoH5cRKiFLPlPCfIS7KfeuiT/Crh4
ixeJPTSbmzGiT+J+KqFe3rRH8LMmw+YVByLTWsA4g1w1JXM6HOqDu2E1EFI069ezjMie2/ErujiV
0KLIJ8Iu90DDuCPXx735ZTz2227T7uVa+UB/XfMRElBm5qaQqoYevyQo5w1fhJTqa9TmEIgULIBJ
9+KSWcb5ECIE1BothsQXQjHbMHgofzY3kKECbQdmpCIQEK9hR/ad06KT3N5gd834ce1eAMeMpwMn
ECIyre4g1e9kMeVwgr1a03gsG3eiTF48AFl3894yAGqxcSulYmapX57hXr1sJ5WumbOExHQWsguk
y5sqw09uzL0qph/KO9KZeEaNSV97/uIxNZwzOib7Rs+/4KsdboKCgVsUSY91tvSuY28YsAR7yD0H
Sx3zxmn/enf4pU1rmoV8A1bi0RTcFtc8P6UXpEbaiQvmIQ1EA0ZxFMn5DYvG4qkjX1eWL/ZUnAlt
KobUzc60jectksZaWLaHnt6PyIGeSKypeH0ePsws3QRmDED2MRS5Lc9EITqkoD+4oIB6rrj4A088
xmRLTNwF8jkHnvvNTyju0Kt75cCKyLN1vY6scUD8mxspLrCGDsiRCrN4aAQn52Tr3mUWfhMajPte
Jo73jOTVtQBatsRwVGT6Gwv/2LhTEthNbectxJWJNuHqwrK7FVvYtpmoHavwJaRefnxVwpAskuF/
CeYgYQzM2WUcmza0v1EtIEas1ougG/6jLglQtQ6V1W7dCIclVq9khZkaYvILKWEOl35PCmDDubrm
fzkoWYc9dQjnnVHOiKhm1mCKDE6RDhfBnoMjsFwxmf+PokFcPWCxUTY31+Y71oFmqaZaSStzKEmU
rury1/6zW7sLREV39j07N9+Y9dgUrb1YOWrQxdpiIByL3mLrf+2GVjE0BoebzofVvtD53LFSHq6f
xvkrM+6mqL1wHTUOeodWK2LyIzA5GbF8lsqydOQiO0t1WLuk3eLSXPdB2dgr/8sU12E20dHDAvdG
Rh4FTraja3H4PWaIyPdNP5JNhhqPt+g/qFry4LvOFVFQ5pZDri9ghU5vdW4zYJLMcdPC8ccTgF7n
2mzN5qo/qm+WiwrwT3JPd/tVeMecfV3lcIyW/8xq/SSZkYU74lnujEiD206l3N/7OMjbPtZs6/rD
pvvfVD+pOynpcSA85zk5Jt6XWaMnncf5k2QNZAO8oCoiibg8OpW9c531YXUaaV4gXwV9uRb+aZf5
20LTXGQZGvp1PD9bFHlxLp1sfCrfNKMPdr4JHSvYslvMedvbQzPOvf83ZmijOKOIGeZAo6OuJlAr
qTZ83IWkMC+xnaSl3q3xvCW/ZkgdlHWMR1/nn6/Ep1JCT6TEuGklnF+PSxq3Ne6Z4LEwset6Fzmh
4KaQ1tDMm3TDlX5GseUaqLFpfH2OdR7h5Mhd75RejyMfUvQMmG+131PzmlSmuqlZFU7frPx3FmjK
6MwkLo0NVMVn5odldayuJSrmFK5KQ49sHqlCwVG9rqWqy3mUVTPv0iOr+GiHSLXkxMU4l0ACwYe4
CqSTubikXCNwqKdqAM1imhmZm9u1kOoy+2hCwjmleEKOfDo+aOVOsuk2rcK8UAzWDoLqJlLn0hSt
UnE4AljTC1j/wIwUsdEqMhbLXvfyW01i3EjNrq/dQUaNtfhuzyGp38WuE6g9yuVLk1djCTx4oIbl
XwfVI6TnJtFvIEOJvyjFNFhnMSnBOKfcrKaTxTpMx+Zx/2DiZ7ULty6bE08bSin2rxT9+h2HWG2X
cGHQiS8yerm7S8N9zgsGDjg2JUE9eCBZ5pGaWPpqBSW5QSUh5cXIu/XWc9DobOCAL17NkIczR1kd
iabrNUOIXpgwddTUzRFzSg7n6J1BRc1YOd4sE1XiVtNgbKlA9JBJJ+N4q9N6s2pN31EF5NqeN3OY
anGnAbbx5TCLDP0dZHDLsPcS76fF04WW9siWRzekInl2JBWnAkZZgdFoxt0XbBpZPMQRnUpd1+jf
rS0jXAH1bwnd07AXrnLO8BPyR0FnZ0j81OC0jw/lqCJE9fOb33Z9v2yiSg5xOYGmhsepYwik8VDM
+tKiOAFVMGgiK21v29nXkRoVCm6lRa/0VUnQmM26bpvgMBh1OhWBJDo/b3cQyUNcmcfCQPJRubLI
YLDpiv0GfJl0AfMFfG2GTKqWg068vDzwmZLGCqDEvOOc3/SWqzcMDeU3B+cCeH+zsGYRYr6lYDgQ
890KjxkiYZvdVYP+F9fQqn+eyi6/sUKx7U5rwAribE7pFAavlVlvZrbTm25VsIMRppAmG4pnFa3t
6/lIit4lcoCmcnOwjzdyGpS6mc3Skn4irgkmJXo4EwP5wN8Dy8F/XT8PwdAhvORcOl5dbOghjO5Y
mxhZ8nPKFv6Ye8DDo79kJectREjuXSZUlM45XSi0KXTfHEPFMfkFtmcV8088YXmr7pHzBeLlx2nF
Ib/RrmsfCt85NcUA3RsBL0DABffPOTecKKVQr2wFeuLhPvPz3jv+LUzLQaj4eM7qF9VoAQGzzKsW
gGVX0C30hBPV7Pt1Vwc4zPn2QWqjmbHk28F6kt6whxloMd1e46bnIa8qn4w0h07u+D5QqiYVTAF/
GAcpibjK/bIVs++R5hocaln/neXGERtRGFlPLMXcT5bPyuRN2SV+6a6SQpSspO4BnYcu4Vc6n67P
MIP1y4b1nNJbcadybjdcBUGRFFa72v1shGthl9Q89kX2dlZMbaNC00JArRRUF38Z2y+1FTm9JUVm
ILsIqkYC9C+UEbX4Xb3SXBTEJYHTNarYCjZJG+1gr0SLVTxSDUiw+U+Ap03KPbGomuoozUd2jbM+
EOKa4xEtwxZdhEtVCvaq1lhbYPu4NeNq1JO7ro2HceufJ1XeGw4atfOlWWept6/ZgDszo+wTkR0b
AllUwW/OiBBrBqYMc5E9yQhS2wjjPoHyFjEh20k3V6XphpKaFaxJES81Lh540hYjNvkXvGruh4Ed
uPYM8FSiY5xUrOr0Em3PWDx1wmD59SaWX6VCvocsmNC5WuEmOzvWUtN1LoME0YVtd/iyKRjoWHq/
CIHlcxqlK/oZwa5y1X4fhBc1kE4D/ggECaOB0uoacSwOQKP40Koo0aZOEyfLbk4ukJ8mf+ZAhtZl
w0DMte84TwoyTiAYQcwN2InWMmuedpZFSnS4q+jvkJ1iciTVCq8FBCUyv6+fmhN4R157DliqaoXV
BsrAywxZ67wgHH8bAHLmnOczV/E2dRv/JqzaKyvGUP/38UsJpx6zSY9DsKCbty907Y8/jLu8yxWt
SkKVtK6dvmnzDRBPeGJCweKhuhrwrleRHdwuAfgemDnjmwdnnh+DDpC1FT4ebHkI0m/FgLmeFBf/
D1ruzIB/R6jh0+OB3z22Y2BR5qpK0EIVeuoorJYRPRrlPuE4Eu0aB4d/9jiHrPOSnNVm1H+RRtIw
TIIxXUPAdizm9VStqaWqgnlarOVu7j99euD62Ld2sOJOusccUW3xzmBOrIWrKRqwj9K9LjUbFZQ6
IekVVP3Fhxwd65NQ5WlMn9KxZEemMWZqSxjKLZ5Tnjq7LJheR8xsrE8Y7F89fJMiaHc1W35hH5Ba
visrklKQHq8n5mRxV9ZKz2gSre4FRNPTb/3L5bcCwWWfMfo5dkhMwgbPcBJsiOgK3+Oi4F4w5mZa
8UF9NDUqkhJo+txgMASHGNaMGbpmyaSEsMUeItKbygf6aqXlaohO5YjgwqAjtlQzWw3zVkH0lg1j
pS5q6YV6J0ce1wHDULTTiwVpaz+wLfeq9ZBtwAd3hQelwNts+ODXP5e5+4Jx14MLxw3Xy73AMLRg
13JxG4ZpVRIy0e7nDlw3a1Ny2cmKqWIPbyx2wqaD0qFvPggv/pkVJZm4lt1z2/3dnBsmzVcG3SD7
lIAA2IX0l4PMIMjv898Y8+BkilTRmxlU4FHfO6txXB8U2WxeM+EHayS4Z+aWrRnn/bVAnmnkiqxW
rppkTUvdub88b0kossa+Yydq1eWnW0s+/BqHwk0nDWQRxVn5EBRG/9bgMBGCF0QGpc9y6mo3otWF
wPMHwk73IoOR9K4VIJngkQViwVTwCQgFvVS8iTHyfqKXELD24O7wx8PI2U4b9+PMmxUXMB6EN5n0
uwJwSL6yBmugd2vaAI+rZPG42ypaZ6PIl30bs31Af6EwREAbx8V6psvcbtzD7htDEYkIp1vCSeXb
72ZaMR1+vwZyuSNkaTqEpW60vKltBK56nW8Cs29AOTG1+E/ltDHNKPkQIMUplcKwDG6h/iaUOVV5
lHH0Zg765p0jJ8HnUvdMDu8B9L7UN5u9UUVWq4GHvMx+HU3EojCXLTHWRn3v112jvahezBm8Bq1C
rolWhe+SbPTEKDWSEwE3CsTPaoLy4LRTCj9S8Xh//e5ibSGpI/GN+DhvgarV3pQLNm3nNgNwM+9w
NCyy+LEpbCVChj/OEgsd5zHXYzMQSGgdyWzhTimkyvzI4MWouyefvhE0PB6tGDEa8WdVbxDC6zDO
Fp36uRv+GSjOVS6XDyV4cf6sz2V5N6k/0FeAXAswsSjS5D2EEq4bUBkx4wkNGR3UBUvuHGmH4ed8
McdpIN8pNVYl+yabV3h4fkGa6I2K60EGOp/GFXIXp/XZR9BNCd3g7qwvlrvHIHhWAL2Dw98L0XzA
rYfw8u+A9EJeRZWNgyOSH79xMibJGnX8rdF6KWn59U9Md4fe1YiWQ0zAqJCQz7JP6voP2nMsMLPw
O1aeRNWLqvpMIL8r5MP+fOIZDzc2ikzPMT36c6TPhW68MkkLcsvXVEHlWdD8559HFPN4BftK+4bO
SPpASCCFbjRZY+CRpa5ycksTEnjNW7JPFlehI+zQ/rW7MxjEstP/ktHK1aD1Hk37jAHiHLvWAAJc
3xSsoEBK+XxKcOMbWLqFrMHZKcPAUOXqOK4C0hU/4NuS210H/PJq1FsKXRAouP51Ffz6mbRAlg+T
x36NeqDzFXZAh8YhARqDY4jaRhjcGSxy1NcxqvCcMh/XjK3us3Sh3ySCvcNkYlumrSTvJssAzaZ/
/ZSk5NQ2iCRtExbu3KhB29KKgKFusi0jCl1rrfo9qHNJgcQJqD7uHpNPg1Zb60dwr5Ko/KTN+3Sl
z1GlDXya30i+a2GzmbwczniX49ysdtZCHGuAbN0k7ZU5iURxwwoV6+oNGopD5khCQagIqcvtxurm
SB1cOq0iksWOWiq5ZBmmh1Sb1nDncXPjhDMbdrTsAGtKCIKcbuBJOScAyn45spBqn0J+lr1ry/JR
9In7wCvRQIDlzTow90rxa+1HMueLmzmqZ7ZPVx45Gnhptfm1flQ6jPeuwGLiJnRPbzn9OKPfy1n5
xgigqhlamqIFE9namfPMcaWAJ12ci7EXAUyFcmKym69hcSALsRJX7TDvNDVNFbZapjoaA3fSWnzm
TkYEy43gtvEMGPR57cdXNYNZJxaTDLUvQR1zUSdFs0H5qjG7QLt9yZ/6qzrDxWMMrimhXepmT+6e
mqE4Jvy2p2Qqp8VljMBTXiPfR+z4EniKymIhUEyEKLJFDBsha+9H3s/WSSy8hIgorLYkgCo0grwa
t4JOExgmMwuDtHpfMJ7ZIMUEzwETUDnLlHUGmG8ONjNI00WIbjF5OXmXgmmC9KBOyTaco+HvSV64
SE0pIoC6dRqa13N/E5aMj+hwWSYW/khTfKMR+BlZogOQUMYgOZn3CCwpLzorqWHujnSvpjAHX2ba
fVX8i5K2ecuszNuBqaW3ivc5E20YU4m0/6sj+rLyKXutM11XK2QRgp7UApDTHJqaeUYLsbdhMcQe
VrsiijYJ7GLpDlzDwijOgRa/opwmG7BGrs26Yvlu9vfvC/rqC+BiFoe2fLiWo9IkZcp++tgyOLKy
50Pf6pRYztHZNHFE9T6B7EdkqMgoDbVBzpDRcX7grUlBYgPw+moVXE4akMmVi4FR1t6kXBrN0vlX
r7yPvHpozxruLCl0qZqoNVpeyic9XZCumO3r6rE0TrLPzqAZAFdjfiUHaY4rn2d0KUeHgbRSqPzP
CRlXHFzwHsdiyFyq7lTwsa6kLBEOzOvWnO3wWzudurGHwGsHi8jZlEECjsL3aDRmeb1OQE+vCdMo
C8ZpqNFHQJpvmgHG++qqnEQy3RAn5qcUZ7hvMSbeQIEQyblXK/oB3hbmIjHYKisKHCN7Or1i0vVb
EC/9bek4lVsa4jFin+38T1DjOy6bx5YCkl6Md8DmG97E8alg45+SkbbQdW4YARoqTL3dIilRQm0Y
7Do15DQCow61lGLAVXvXsxEqktXt9CnYuYI7kzsMvCq0F0c7A6jGruJnkmGGKvljs2YRLK58GxhV
XtLxby/ugT0m3X3+ByYgIhUdbzC9526W+yk+f3+av9Vo+fooZzmusj4LnHAw2gG2KOX7OXgV3JJv
irPLvZLOOXxX0MMRfdRsVgj9XZ/eXiqej9Dn7iXPAgK/kusjfXPgGvqCn5TWf8HRu+1GfDGmDLYU
QofcFEokEoWXRdEXBXvY997/b84T4tawTedYSK4Jab833ZDITCjIj4RWa8MzkQMt3wF8AgDsGSpd
OyGk2F1fQseuvpbC9Gfz34BfNl1F3XweelPv6pNIXVfs8ByMSDm6J+ds772l6o7iu9M5PUWYzNOW
ODDZDI+IJkNk0Hoq/T9VftY+A1oH3x2ik7McGeWLPIYUJjmB3ExMb98pX/3VAKd2LM7vKaEz9ijw
QGRvmzUdGVD0y+X+spiQw5Xsb9Fo/RGs9dDnIdWbESvcuEJjyFO2MK+GQOp33yt0UCnbrNduVso2
karYgvtgdlCu2mwkzBoUAsSpAD7eRTjpvABv0khRYRBY+3LyBu0dZwf2BhL+BTWuDTmFMpaSKZmC
5XKtH8BsA42OKxMmube0cFjIm8WcG8Yek0spaE/8ie/7NqJgSPJdyVpS16L5obClDYQWNDGGXXvy
ZDW/HMBeJdvHFhX5ZJ2ilRBJ6pPrg8WhWSkacJd+ykYwbMn14N2VgxoQncDRx0eH362irlLkBgQu
QkCk9tdRS1hEWPIIVgmGdb19zcVun5NxmcHVjq9jaNSWSt9K6kGOTcCjw5AGD6SGULxn0bOQqH/o
7AG6xw6v34wY3UJwbv1OX1GcnXx6A3bGTrAIsijM6Mkk3U3YV6+9u54uoDeWxRGAStbLtdAGLoX/
c7tT6eXcFRF1mOPLQjPH0qNwCJh3ImBdksSZ7I48J9JVfun0jgnWftmyXQ8CAMbUu2L+gQRE+s5L
E3WmaYtRnq/LwoHniSzKo68KbAsWHKl78Tl9G19i8e/Mvc7QXfP8rJFFqM63g0mVEH+gmG4j0Y3l
3jo5j5XPlKU2yGhTmZqvCFvhf3qJXt6/p3nESvZTBUP9hN8f8ov10m/QyjvAWHmeoWj2/o0P/r1c
6Fp2o8eAgrnYbrWqRZ6zNj9t6narNPP4/WrNGxC7Mk8vRaga80VfHslqpNjcXIpovvyaehzgyFph
F2QOwPFcR5neCuefcCrjPOZazs+nkHrl6wwJClWBptoqvoTMA5BscvvuhirX0yKJ5s+2HsM4ml5f
+E933tRfSZ8xt7R8UVbDhBInNoqqtKs6gOozn2cGGCTiKNcaKkls2Y5c9k2fFIs/ifwB+7p6MIy5
Z6M2m3cPDBI9xbRR95WQxDwCddXvKGQgMSo9flBtbqK1poX55RAQvSOfg66XB916EBJfje6+HpHx
gXmMKrGUH6gtUrjbFM6q3bO7unEz7sUB9DpaKZymwbVWZ7tgA1HsY9WugJPcHietOQ3xFa5yIefx
ZHHLUZBm0eHT1V71CidWilMnYWv4Kbhvvt6adAJZOYG2F5iQkG2XOgSSpZ7hXpX46U1Jm7O1i+l4
wIQQ1aCkPTkfFPQpmdzFwB5qmKVxvvLE+xbnH4BQM14e+JcGJCtpL5McDMs4GA0E6eGSW2cRvpiS
yA7Frqqrfz0kVuxOYLdbnijxe2tIjmA3B5vR00vKU1LfNuY36MzUx3A4HEw1jF091hjwqfuy24ao
NuXihbehtkAIp6FcJCF6AT3soLBVJngRVUhVyK76hbDNoc2OViZQMkUS9Ejge47jVGDOXOc5fEpi
M0qTbLnG57srvCWK4D3GUF7qEZ3p1w/IH3za3uzg9ACoKP8AT1vVpAFggyAtg6SZzf+C08RZV0F9
6bk61hi6gARJQnJMTXpIFFPNrqD2OByvZsX1AQFxj+gBIDSacDjp+uETy614xAcbfLssXXOEHugP
WRG+7cb+2oHm1foPNm0MktdDKPuc2sSoq2s9d3yVOcd0UbshFIzsG7AO40DOv7sDTzPmP7ixb2Y5
RshwVHrbkO0jVbWBE+baLts3lLaClgSxan2pNKaAAu9piNq3Z3UQC0PPBRRkJGdS+M0FDf0ymy1R
Yetfzldqja4OZ3cOj0LAQyknNdVyrhkp6WbFUxP5RvnaaQb0vC11aQ+IE29NWzd8sy6tR77T6TGi
DoX5hA8B7Rg+tpbbuAUWhajbWRBEFg2yNw8pNMAMQ51n2JnbU/357ZsNI9MU3VdCwLm+bAOH/76S
Dfz07FMQUjJhzh2x+usnGhskin0wTLLNgPnvVMmQLUTqcebeNnjz5hTNZ3XKi5VSQpq6pMITE0Tr
cxOwR9THk0LaFNHUnIbXhYQPfftKvhoXSYqnJg+e6PYmRTGLKCZ5vQYRmHQrSx94CTavQGlijG6i
Z1U+P3f3fgeP0fufV5XQ8OAAWr1bGe6Ms0PFZ3r9/RRtrQDlJkQ7zuXf5vYTrowwFGynbAU40t9A
7lHPD5pcu5Q7t0LRLx8ruZXQ7YVN/GDAf88ZthSao8jP+qbc+aY3oNz+XAhnE9s6WalPV4IBR3P9
1sbdTb9uOtEW7TGGj3VIXwO/J3brres919BYzF7VsA6sJ7uxEAijW9NrHn6kg1MU3xwQAA0xstpO
dXVFJR3mCq2yBrx7WPDTFxcrIjdxryjq9TVHi2sl71wRb9bn1UsyemMu31A4tOgG638skR1s98lk
k3Il+rmLSLyP+T3fU4haEY9JQIWBPIB5eRn/cGjJIV6pukDClu83LqsLbLZ0axi1ZqwxMX2/nWKR
fVEHibety/dzBxRGKrhFRZiuPM/Jx8vv/7rnKMmkvbI8Qirh7c8sDiVIHMouz6itAzf4vQEhX23i
Uj/h6sV9e9EJ/lVMxnoYDHkd33YUbN6PuGtA4SM0Ey7V6eGUnvxWTOogSHACCMktdPa5CY6qwKOE
iPnCIFP1GO6uGs03+96dVFWkkWeJNiriDSrCkcukjaBhw1U84Z+egXAdmMxEyJ3p1N5JcKTB2/MY
tzhYVjGGyMhgyOqnuQULbvNHuid1S0S6lxaMUYe9/HEjfESAKBlUvSRtPrOwXDI0AGlaV90oc4JO
8Sq4qk9SHVBrTamEdADcrBDiuqwmljPoZ9ONQ71LNijGGtCJR1aHGCGIopzGepax+bQVPg1HQAf4
W3HqbANs7WlrODJYzQu1w2G9Txm6J+2MGCMTVul1HjMPsWC4CHuOPEpETYbXhQ5cNSJbTtKDhdtC
lLBWTgvSJ8d8BF/H075sJED26laoVMpx4DtORrUINpngP2Dw/0u0ejPRqRZaLlJVnx9pvLGBhevq
1kQ5s5/QNnIBnZfO25XP2eGV+s59kHIYUsmqkq+DRKdAE3smxEwkcFIz9nUPxeddVEDb7p9vHrwa
J0rFfgIPAW2GnCyVyUqV5bHvako5e3F4sgKd7/fBGUc6czwOBZMvlyN79/MUJj4vWI+qfyL1hI+b
UD5kSVwNY7RsLFG+YJxWMzewy/aAfAvarjNRousbvztxAItbhmDHDjRI4YZ1ywn7vUqQIZ+/QIaT
YQpkVXHeppTu4ckFeb39ok/BjZRG9Z2wdJ1tQ+oxzCJahu2AGrrqRC4GrDlfQLoa91MrFN0Lnzw5
M6Kcu88XNf/YOr1bE2/ivVjUrmqViz3KBUnDOs019Mz+coM5m9CfvXPZa0sT3yC0eJO0so5yfJ0P
pDuDZN5iMuJyjwnDz8bm+XdUD7x4tZEtphfAzgPyjAlWQMxewIeh1ryfWcFDVMK7ll1MqOgd5ijC
HNFMLy8U4dMJjwSlx9VjETrTZoDD4DUhNWQgbzeIVDx5yJJLzqRTgTclMmOquteqp1gtCty12b9H
kXB/42Nn4WYBbnQ4F+rMtP+0AHBHbGqTu4Y5qI9Fm0xXjipAxwW+Sf06pVwnTuXD/SaMKjwRzJ1Y
jgBn7BO6SOnwBcpLAiwyNzjKlLtw1hQNVscz7qfiVIsS0JV9N9kSo38aJV3hnssFnPUUwEZXSVvD
Iw537Ar1GktBh/KabH48tETvqQaovUV6DmpL0uy2HSvOZfAj6g2uVip/FVxiAVvaMvBzZrs1lOCM
Bh7nKJrYhGZhH0oTrj4HNWH5J3P3Z7yHz8t6FnbCYHz+QJDfQ9KaLzVJ+nZjN3BX4N9zN/kup+W/
cJBhWhHPsRkQBc4b3jvyBHhHYJGCy7hr5W1JYGrQ6TeN78dJfLM4CTE5lBWmSu5kksVnyDSAxzF9
e5x5Ewn9fQh80kx8I/Jkh+1xacio5GIVkVa7XD9+GnePHZCh2bBvS7Xxw3pB5l/+FJbFqo2f+Jrv
yIayteBtvf48IDdmDLBd80ZOzw0faIkHW/egpTSCTCSPybV3PDzvZSm/x2SoWl0qnPI3CFx33mqM
kf5Oq83r5CXhh8E46hFlwhNqndRTfdkRVmarlmf1u0lrtCTRAGf4zytFxqtLjfOAI4XkFt8z1x4k
iFRGzqeTLGIQ+gGqew/tE5Gwq4S1jIl2nj9ZSJ5RDzYsSlmObKYXW0XwoUgN2b6iuQdgTXt7gStS
BwN64v1cBW4CDGQLhvV+jW0dPnW3XOREsiePMDCans/RZ8FFiEecK5dCkiz63g2RH278ikRDtcKU
bhAW3BWi2Dijfts210t/nvELnpa1J9uH1YGJsgdXJ20AIKVo4+fa5W4JKWaT0169CETUPJHkaCJX
pvAZ6zJXZjYycEMIaRW/rkOZDn17We29lVfwxt4n32Ow+XVOsTAwe45SopZ6y1jDNSBlPH0/SiiP
lX1tLG1gnPhZE7MtPNVaoramMkfO6swxNG4FOiGlvCG9YLQ4xrTzKiNXwbtHFc4d+c4WKX4dIRiC
6cxwNJcxVAz52UpZqdU3WR4orD1K2Z1JFRJbx2J18H9A2LMKMTizgXdkG5Lan45iLGl4BrkUyi5t
gFZ2MQLt4cPVaSAxxyC5vUupf8WmnbnZl8WDU9OIeHHCxVGVPIqHpz6jj1Aaw4ju/+5HVT1wz4Zv
Jdszs0nC59VNcYOzpYWOwLSsFpRdDiIaaGy3F5klCWRXxwxkjrTSYzutgTE9r8SmkngXUv2CDtyv
Zxbp/ABMMxXKGswJpLN0NSBbrPzriCnLGTADoToeidIc7idGctqcvPv9yQYVxEkH96dwj/gTVvur
/N7uRNIcNuFqj5vz/amLNVmENHkBcbaViRBUotIhZe/mF09KZsA+mzC8HQDK6He3fecwciUvOPvE
mFo58k9LTzKIAg0+oG1DxldExfXxkEv/6t4uIf93zYusJfl0ow85VYJXAFJcKHvUbk0MThixy51a
hh28I/yZC6E+FfAcvUhQZoIgiWGdVm3LeEqu/i1ERHHzyZMMic4ziwTBr0Q0vkG737LmsyyblK7d
dk6Bsc07xqlOyXm4JDvs6r0QanzdlZPxFM2BDHd8ZJOGfxjWmTN3ljGD5sPO98dAuHQHXfoOGIL+
mSgAZ4hddfj+hhyvibrivPzyCleZcVpZf+UQSig6ReCI/p6DPkMOBVQ3TpQ8OxCl34AV4/fX+8po
M6YcNkEzAjB1Tw0rPRl2w9OtkUfpvZaPe2h2rMT/9G9wzuecioeh0mrZaAD4TtruNxX+bS00B/w9
R/cpJZxUIVNuTEEM5mphc+/ig670Dmd3L3hk+5uZ0hnwXxrvrlMLgr2KAkLnaJe49uBk4cJYheU8
9Ej1R6FWndvQNEmHBdwOf9FVq6AHSZ808QPnZIhsHL5bBWvl5zyKM5iIKuj/3oOOUJEIhDzAsgzv
VKk6U5kXC6HOOCNwALWGvJVrpbVO0VFMlLXISSAukGXAgo2iMgucIFBWDh+O+a9l4acOopfNIwGL
Y8BeV8KyL9/MM8eFgugmQX6rrEEb0sXbTlYnZScVWZnaY1G8srWCgImX9HQ6vjCUOA1Xs19IC5U6
W/ZMdw7Pi8fsu7kmgsMyftfjmUKkXlxYEnq3n4e/FrrgAXL3JYZvM+lOVrrZ6lJhqUJelvWlnglo
z/upXV/MPF4jP2AIhJcEm9Qg1a/+OfenO4CuLTFtEM7Ilkgu5mvPkt7mMDj38eGk0SfI40zHvqNR
5GeCV7rjpA8mm9/0G5EQFscZTJCcQ5jWMOQJZRJlC/11d4xWdnP6VvbQezlY/Ne7hpIX+6qYjPZv
TIrPVZ2goS+fnHzzup8vTF7LDJqH8s5aZOxtwjUp0Cgno3+0BvlS1sOtupSmWiD+egNv+N9O0Ykt
bEXw6G+09VBj3UXTSrVIVz6MeYtgdprR0+rJnPlX27SYEhXoeSLm5aO2J6fiNFlc2LElb1qP1SAP
5d3+US8/M9WZOgNz5dBkW1UCbtsdAFOH9y+hNoCg0YPdVn18qfZSusaum+ZMZRhCPi4Fl6ejS+F8
KFDRZK1cqkb0ekvPoamC1VCc+6AoXgkQwQYCepORgx5RPd3UA9dB7CK/3U+J/9H0KjTF0561qG1d
O+UyDy1/pylhhq+eKkrYrJukTl18wsttsA1yQdSfvw/KJTk+OLerlyT4vqNbBvE6jBAOez4vE2c3
SMTY6y+PLKRznYTmcEaBq21ML0JhbUnrbq2bV3NgfoWaopCV1w5EBOOYYhbUsPGcnKV+5kiyvNJW
KHx12zcBPcywY/JsB4KqtxlvQDWSWUGxz5+JiT1+pZyheu4/3i7PRIVr8RnAcTFAuLF0onZGX8wY
KnPWFzQYGnUYGJaAuh70CFIsPh0NfCXE5lu6+88XAWC7L/W38I8ebKb+PocAQ5uXU+ZNvtQWSKEF
i6pJDFUnzbfbMP5GL4oKkd5XvTaC+kSxk1UMq2RCl1BG3ASw/juicod5EyqfW+/2AGl+acLFGIUO
88Yko03vsuuF5+PolvuY/YKlHr08y2vKdVBG99FHaxJ50ibhnIk5tWOJy8IHYaQUFf6ptRxHLNWH
Vga9eZgwIy2wMuDXk91Tp7gRS40xpI7jbnlZP8eCMz+n7gCp63zvMR3Xn1r9sB7WfOQTlW504po9
YSUJY2YwuALhmkvBpDirpxID4ubdIoEmI8VcmvIpbOGTNZaEODQGJBiKJDC/tq+/sLHonnz+5QZY
3saRH8eGMluuOTo4di5q4lKInu8AU+Oqd1OUYf+iBnduMEwc+ADDQ3XHRCui/83cUmmmjTyI21aQ
sDhlbnaWKh2oEXF8Gqm7NIaIIKMFjZ+2DGUNiTJfQU1ueBn5gp2Wo6M0Yo4Fu1k/NMBKE6/yKWCy
3rN6eHWyLChgjfHlG6lSXqJdVup3izWoMGSvy5SnqxieiPHbsPbHIRNOX1ZvmOgViqmsi7m6VsoI
9Tq5LQq4gK4iwuvPotPNxMGwKxlEsSWALsiQvlBfdQe/SrvnFC3NxtkX0YXW5n4XqgQsabH2X8E2
aspaCwjB8ZzT8fc38ZMdLOJBNznKyUAGa/5q0OfLOwiTbsbnBbw8S88mg/0j0eotv9VJMBIPNMLB
zdNtR7Xv+/+Ffwc4szzw4KSowfoatf30Ibs8LAa+n4JF/ydtF/M8eNHZhOvPimPkn96UpOOkbNG5
BWzKV8glw0q/34/5ekBd/wFpA5xYvQ3wGlsNitBtORowzScsTqvHUifnKYYqhkDDVAPdnZ5mnOmj
13o+lX5LKYKZNinI/k2ximEOweDOdijC7SM7BVjxRSW2oq8MEMTLNFs+AHyLJYDRkcLBIFNonfBU
UsD30q/eE/EVUrf6R9RayefFWPDGHIcRPXegWaiS5XY4LlY1w+h/d1urV5dkts/OEDwCuuT0JCyO
aB70AckeAAytcq8UTZ0H8UADyaiQzXXPe81o0KM3bdNopnI5zgHcIkkTgTzXzi0eToHQmF9TCLLZ
kZ6b71fg0EJcrAS/w4nhP2bo9LHUaCIOkR0d76yYeFp35VVZ3HtSzKsXlf/95BODpaUQUxUyXzEx
EaHQ6fuLwxoqT8WdN2viV+v3/abByOhmaDwLs2UCDMOXLDZ0GCYggMnx4npT7WA8KGtAakUruK9b
Her79FkFb1GkW21bq9hU04w1QIY+/gSnlnVL/6mJ3TB4bNBWjpOVKa9C18Z3BglSvCszaldSesRg
dtYQ29ScyWVIvD2VmbnHNPMDtCdI0x/vmz91zCVTLm2CY7su+BrS+qY5Ia77MNKHebokFN4C9aNy
SRJHp27eERtib56fkPaEPBipXzosP5ub3RXbWQHocdz42JbTLUQj6HGORESJvCwWEdDNS7eF500U
edEC9SmLOdHtxB0MrHG8n86gRqY///2foRqaowdZAebvMvnvUrf6KZQFAGL9/EJmR6tOkhm8pL/W
WSSy03HziofZzf/18n2rL28TsLem9jxqVJfc9m6oLf31fF4JevERUUvGH9KW0Kqb/wBUq8+HbfYt
GKzwPr0+uezlvh8QKnULJrhGwXGviijVFwqSzjwDkLDEGw7dfqmb20fnj9l010MvapH/r6tTzLo4
3xhoiUuqE7mGeb1Qol9DzbOiYtBM2pURnXzK3FMX6DTaWiN6kmvOARPTzx9JWjvhSX6TqAREjZZM
fI0b+FZ6A/JmiTC+ELwX7TKTaShNnzmmJle63DnARbQ1aEgaegTJrdtQAUp8sF/aEdIC2bKHo4f9
5jLGEaNS3Iqz6KnhR0FY7Ug0D+q7RXUqJZYbH1AMYpbuvri4216U9s+OOjKkz6E6B4bi+m02S0Jr
WdAX+buZQGaTKwxXa47s1No8nw0tG7Jc++yB1U4YX4vowtLB1BFzMJ6MFULMYnPytKAZpqGq8/Op
15N/7FSYCFJMwWRGwgrf/gLtN2I7qS/GD0bj3ikU0HWXsnQOcWAwLGNKi86ox1OBS066e/VUewqy
xvWSNi92gnHICAPmONjLkPsPjTEUVsc7NuVbh2dxQXUmbs8NAeciu6sHVfEkLmuDlH7b+BC3cWDG
g4Mc4q3Kx4hRDpSWRn8aQDuhYFjb3gURWsYcyIut/gvXrmrHgvYJqmfuUvOgUisClxwkESZaVeiS
U0WZZ683mawP265r8cwwpfNkoW4au2BA8mvBYvCZilQuWyAJNBQ7J+XKGFJCwVndNILUAniiiduq
0V0k/gcS6sYRHwb6sL8AYZ6tiYHj3go9RogsiJPonPPKP0DAyNojFVAnEmtu+7z2927W6HWqO1LZ
gVI1XnCixSpx9FgHG58f876ypcR7vYb+92J0+NmkaseIc0fVrsJ+g1YgcgT0ylk4bD+clTGgM+Yi
VC1yIa23p8HygSIKV5C1pG3aQxGHNk1PBPn5lOk/nlS7HCm4R0SW/Tng/oU74JO8Ry6XUuCbFiVy
OVYOoHjUzW5rBTVCn7E4iusZApFaOLK+lSS6+0ErExHJK0afL5PIoKJ/QwMDITJbVA81OHy1UdsG
j8LBPtAJ1BjPe521t8YohCRon4qYNo3v3T7wGejF8Qa0cMsRm8Uag3jummRfdZ2borZzOz/ieUqD
atG43loByEUT0K36OGhaLlzAxXNTZD9PuVWHrkHYHX8NLXqeKe/qQBkGZCvFNfbmx5VDkQyLuAHv
QJpUsWCsJWlEmkLuRxiIDyAFtkoWDPqLFfk8Xe1c3a6nuxmNARFeHHKGLcSS4gC3E0D/lMTHsoLC
hSVeTQ5ROSk3vOvRclRnFdqN136O9ejBG4WhsiWOyR8l+VAllXyPjRFomVxb8RDFbiANPPcC850A
bc8HE0C6kBPEwHngGI4upbGKKO3CVwV8T2UgzXJow5U6197ma4cMlTkbwwghRmXmxy2o1q3M5ENL
ivczZphKfMwcMCQ+D2W2ExBeiOAnGJkwKO4UMABBRi9acDCyYpDFI9DuGPsu+0Uhd2qlk3nWDPEU
9nqXndhLmRx7FIqT4tmew/ANhOGsQmtOs555VftZLFBCzU6HVQr3ZZ/oSYIGvQXtTIRHruuZRAvd
7+0kX/rWICRB1nR+v4Yhl5tqgPg1QCW9gJE//XEIzblfiIEkwu2IZfvlCJ2xwDR5Pqn+odAgo+h4
kDsM+JywIhXzJPdcpXSysyj2T/HqLqXER7KSojvpY5YHWqHPvnfmhhEUrfJIyMJywSMzbjAAJqbz
ezBDdWW+3RJLt4O2QWtQkGYvP3JvjUJljeok57jmzjWw/KENY71N51LffJ+s6IsIF0lEbLJ+37fh
67xM1PqnjPXFGYDvvLfWrF3Yv3YNI5HFNiTFHwinJBMZx/TJL0RAHBWQCOeBQSCwqzsV0PrfB/2k
7KGAnp07Rp68Hx0kImU5O66QifUjNHMm2iHt2r1CSv3zVSMnaqRljprYWgGEJgfnQdp8XhqMeIN9
pNsWvHTaa8w/S1WVFiCLxnz9iiCjwgR43/H/eM1MbSwK973EUDoSCuH0KSu89KvkVIKq4CKrJyL8
XrFtuoXeG9Z8v+BfV6qsd0900ikuqafMZtMy7LxGLbEZyHzO7ktzveaaoDtjldShnSin3ApviH7M
fGpvr2OUzth8o4k8wtDw9fCwxoor2Q9aEixhhlZfmOXfT0Qh7kcBCx6ZU1BzHTRP/jprX/+tyuBJ
FETgZgIg5pUpdi7Igk+7TRe7BQDuOqCDYfyt4MexgZ94SVYUGBmptyyWYxge94NH/JoGY7/8DjxM
uZGb0UvRuzuv0BwqraOFvQmj1jGoMAHIupLUj0gKB1QE4wmhGJ7vjb+zYZBRFfJg/94grNPuYQwj
97pBVLZUpfN/P68CUpbnCZSIRaYG8O23YM31C+UnIQmHAxgHun9/dhFG3u7AL2pdZ/V3BkzmPKBI
wWh7Lx8TMzTmaS+7nzWdJIt05Y4jlAXTtSRC4qLql/VwKSbeyKWEHEOyCPxjAET/wD1Lg570YKIp
OWampUowQvcjKJiJB2nB+dzYIaYhAnV4sY9zDeuX5adgbCsGtUTEYe4Xv59Q3gwBwS4rz8wuxzRN
102nv7arVqC+FQsPgayokRMSjLeOphxwuogq9wFgta1n18+8RjJ2ho5EbopveB2o+dpdDRezAWHY
rBz3DximPfjCj83hXuTcisdg441OI/SUTbfW5w9wrHw1qDxAmbQFqaJAoFV4qedehtGajMXxw8Su
FtqJW5Yvk/jYwCl/C5elFx/dLldXcbVl56XoeRSlgKlzPy8Nn9oF42FA2xdkEvkI99TUjd8cLVbL
+aL1S2ADHOBEwxky9dO9BQJZ8sgzjiDrTJ5pHrqaXydT5e+ZyOY+hGhWx+q+4eRfjRtGMbk+oNGJ
9kFD3sURxLzk8OYsvSP/RuVEhLGuGFykyENC41VL66o6ThsXEmz/zn0wNet8P1cR4xC+X7AP3I96
AB1p7QTa7o2saatyB+v6voapYegsHd9JzNrh+pQgT+wPhJz8j2pN5kBhps9QmNp8uRp3C8IhAes4
Jm5v/oaIfcac/6w7JLz6YhcBVsaHtEYYgxMYhcop4GVP5xiGhKuB81q6T+jH4zpR0fJnNpWXgX56
MQ7X82uWjIZkOEvf3AqrnrYxsI2EgOIlO4/Rauf6RfC3QJayMF7uLSQJHjDxf2/7r9hpl1B/m0tS
oR6u8OW/kenWlP4HObxxJFnUBJ+bsm6cHj6UIFlwKpgCqHHMyzO5wyxwEsp7ozT+2ELXIkdPtz1y
oGpko/Yf1eRFHqSxwZgfiLoaA53dRS8pLKEwM+KspDcMp9eHWPEFjW9J3aERN79T82IeVQ+nPfVJ
Vzup5+L5KzRabHYiDnojS7NUUDvxM/091gOCdIoTqAXCJJzU08VGLZ4bc1EhQOvSlEeduXGBCEjf
jwi13RYyvhNXIq6kQtg/EC8SpIuHiolIUX6io75J+WCYaD36V5MWi4paoKOrA+AamYBWuTeLbsgg
X1WT89okwI7B3oEP9GPIhcJWWjPLcsvroUICbMFfM+QPWbGzAVpeq2F6FU4QNimdeC2RebwMuyfK
4SATOjfcJRpxFIZ0ZZvHuFcPU1n+3ajKaQLc6hbPQDyyOeCfqIgAm17xDG/hr37hqJmhuBn4avqx
mzFM7YmDtUWYTSLRp50Sz+ElJIjzT+PA/w9De7lXQKLKw1jLe6xiUM/9z9XihU0XzXhelZVcbmYd
2LhtYvz1pio6GOvjcz7DwsZKadLhYTMov2Y+xs2KTuAaq6Ho1jACFeOVLb1aZHhmtgDCx/fmH7De
l+GoQqkAnixmJexQrNe1x9/e0VXSU0fv8T66wmL/j3GdvXWku51ESiu+9Xg0HZ42di5rgW4KCjxb
mQhK9l9D8OPpSpA4MVDR2wPTle5cO4kjz7K0/x8kcaVDD3WZ/BINFAVxODAKmiiMTdx0QvOQHWvM
mKWvVCxDNlBXFb2VUb0OLq9OS7UiYqTIKwwOAUQGYoW5jTZe3FeBnSSLrju3VB5PSvJ474GslYYf
69Ryv2p7524KSA4prdw2JxQq0ng9jlnInBiKnSn3YXiNx8E/M7g0rlgjY8OMeksd6Is+3ul3Ft2V
edas3++nTL+JiBKBsK1MqNwUuKHHwM3bahTg18TL2jzNq2Ac1qMFwJ3+jwz90R+/eatBqFO4l3HZ
ZIkFYbSsfPfUlk4c3lw+lKq1CZLEh+DT1j3GHI/PHBc97rGpvtvysnpdja74dihBk9IZ0ua4jLq6
hMfy67IjfgDfeuNGKCgo+xDNvCfRN9M71cqxsL0p0dvYAcoaA3+7mWkxK09O+GDDEiE3pNQOe+as
JHIG4fonnbzYSeZg+xeoGBCaVUbYzVeOw5UIUq8vpvw4b1QcIeJYTN8XLjab1IWnperCFGNSx4/L
XLhO43CP+xn2M1Eodv0/iNBBFLc3co5MC55RhD7EZFnOAFG1v5J9nECTTXTN+btUz8WCOywm4UtR
Jxrw7cLE40ItJwDR8iusRrNjIVKLyP2B4DllTFcix5lRYiMg22UBxDmAQTEnUBXFKObKZZ16LDP2
mITop0bTIqCIVIStBdWjdM4OnjGpeHIdxXc+Q+D9gIplo75pmbok7twfBDpy2Up+jgcQBuW5xTJJ
rI9w5PMFWQzb7Lh8/ecCvQt6EcWwoKXOEmoN/ANikDf2iZcCgTCSwwiE3uSwkPSsiR0T6UbXNhe9
95NkRlPs6rF8I10OxUjKoF3cN9EFL+AgubtVF1ICAhmbIGio1lfkX/CMgUD5OboSqra2d5zZHaG3
X1HaJLZU4Gq9adjb/mycMd7dkVmzpTe/l+bs6lPrYvYiX1/kQxDGW8XO0yHBSWLyJjCIbyXj3aOo
IAMgVNLmzt6cQ0oB/S4qeqJYaPC7c2QUF//L1vJqJghGaD7sunrPgHzCh0jlcHWBxwT8DCYoW5RX
RY3s+F5fWDP6YvtCp7tr/lkLZZHvRvU4KUaxwHgG5facyWkvqoZuk7K6+2UjuII4L7P/qFH+pNZs
dwynhhALi4i+iVgOKovTeoWfqpLkk9ItJBFJ/ZfrT0hmd+gVVyf5HBgN90qxLiQ7URNuP5hyRKat
LI/0l/YXEHTZZw3WBKZ7JpHHEmMTVkcWOmGTi6ZH+5tcrhJlv0tNQJXvcIsggV3OozSeu+ny6kNk
NRPmi+EQZrdwNtkvn+DtQTCFnI+QQoKcKj4jGpBkoL6Pu3lMTCCnFjlntT71/R2FEJ3VjZZbOTDx
d+ysDWFNOIP4EX0gO6rCV/OP6IXA44+ZJSGNB3DPcc7Hg/ejr2Z1BOS5UGmEMlV87yAMzkVyrBmm
mYAK2OpWBJM8X1y1+RZGqYSw1T0yTkKp9s6fCS6Kef0dknCbv+dgnG7xmezq1BHLSJDxELSTOkg7
drfPfWJDqsztHx1n7MpYNa3Lrhzmh1jqdCw35vyfULmSd/cO14MdCa3EqHTB2e4aVCtsCNclqVlf
SudO/n+ZBB0e6ouMXMKfSogi+72fk0P2fl/9SWUYd8QQJkCDzJyYQIvjtt0pDDojW6b0/sma9XuO
5JkPEwoR60uRaZ06bAXH3CY5QnyLRFiCrqX2rf1M+Js+92RncC0ZX+dIFnYZ79t7O22ttM2OLpSq
eCcpFYwQHDY7G/+qiyPgSE20NbNWRftqkbv+yL/5UDeX0ogcU+rcMSULr1ibLpPQulvEwVkH+gMh
u3T0rHH72mIfls16MCrqr0cKKsHkMt9WAPSjYLIofL96qW1ScZ4tmSegbPOuj1iimQSahFktiTiJ
FyLhmrTwBrHORzYefZMSq10k92/gkPV3W6Migb8BBHPsavzZLR68hD5GqMu1jOqAXqvNy01JaoNi
FhJuKb+G1CvnGxnVL7BEW1vhGgymZDVQL3elm/ZWIoilCpqkllmx5FClkvEUOqNH0+pvphMuFaF5
n5I4awrns+seJd+pAYewP0pyjB5vw5od3FWZR1zgIoeAov3PlgugeX96dFYAtsbwUicL6/ntCIzJ
WfldAwmTwx+T7hzQIXsl9kzww0j8pSl9J3SWfpnqJWgZUm9NH6q1HyoFtJ7+ai/fGcz7mHoxp2tY
x1O6x5syhT47eLgYDZhGQGkwP0d4uCEi//5mpW5JKNIOjrpibFGfUuj9yi9N17ssiIMX37ZlFj/p
1fP2KV4EhaM9nQwoN3frZruhC/xYVIt3m9Tq4EvpsmaJG2pQng/b6GY9aVv1MIXNM6OJ1ZBLqAkw
sl7+7D53tHxEEC5GNsmeOcrK97tUJ+ScV4KIfUd0ur4MCj/K9Nlf/VA5t7vKTKKcmLkv5Ie+naAJ
Fg195qc6jWWB5WAQMgFkhxPN9OsOQnrdFbH/eCrtpESaGEM/mDhxNjeMTo6WV4ppB3tlkoifO8XV
jbt3BiJfRUG4qVfmSa6bOuVn+kvoQ3Ux22BRIWqmChQszbsTN4lcsqFKW7C4lIlG6U+ywzCd1/7Q
VBQ0oIKM3ZhaeG7Roh1DdXWlwkaGIEiFhPbsxpFLfL9QhLxmOH8uo+xKGbRQfvROBy50UUICri35
QNwrYXgD8Kg4F3jTSL0h2gdTOJZnUQuU+59CF32LIeInLh0XPgQNPhRdcf4/WiQRfsJDY5W+Dd35
CreQoAR29Bq6NCS6GjY0i9TKSCcIGQ4L1SsoiJWpNm0059HxYrUPEr82uLOMUlq9vJ7eCfP89z+z
fapmip6drxsxXqw1MstE7sHtbN1STsTP2jC0ZCn/ZKKp314G2OL6NB+CmGDD2ABx+Eb2j2X0kvzl
H7vPhVeYMf+EtUgSvaXrsg+nAXcqbOmaatTAcTTdJskdSaWou47BEV/xoL6EyZOK4tKaJIuCJtcz
I8RHKl64JM9Noyi3kvjiKDNI1k3+7G8JKohbWd+V+a6cwZ6NVqbizCLJaro8+5LckJQALUubBGdY
rt/S+aUtqaaeTIzM0WkMLv+B6JWM/VouwJ/T8x1k+oVmFcGpJOi2fWmd/+M7bU+O8iludK189yn7
w6/97tWbjNcgIEYTd9bcR5jHK7TMuz7iM5u5krHR4qkwKGf6TD4WwxnXECAAbxWA22P56qkfrF7P
6H1BPz9zFMuL9A1tbXb7HD5C9iaueMfdGlXsJLT6N2B4g3Q/7A4UAvqPwUr58fMZ8gwVoMaCXr1E
+3dycr/VHxy/6aqbrY+ohQMj2G4BGLZdpqDhimkXkMbDuL5Av468u1Uh2v37QDuoGrfu7pLaAZKh
goe0NYort9XitCbBQPL8oWNM7bDZhMdzgDlHL1iKh2OfIAoEA+WUn+lBd9iTH6MWR0W/WZoVdJEy
bWG8eJurSNSMDczw2Fbsej/F+u9pAF+vVl41i+UAEseHixi3xaNPIMPJ4VFYcaJC/G7VHKz9TCKj
FibOE/5jx1ivxoPnMpTxyaCwwfZWt2tL9HIrE9xfVPiFYhNu6tMLWbDcu+VRSoPUYVwCafv8BeuY
0+9yE3nbpBudon9X/FnITZSBpRHm7aGDpXsT5ez7dvkvEbornFjd4ka70HT7NI4AleD6bTesNyp2
Hu0aErzrT+AaISreo1sxThUKWByiqAHL6/QH4v5TzqaQVlswIGBh0VIf+GooTAPuam7UDrluLJnM
tRMV+flKzkExetu5Qrqxs/cDCkh0QNckw25c5gQoo45df6PM1+F1NGqwnENOiihkoiaWjwnUsr6P
2GP2pwsSOqdaZRV8yjsC7eNzAYgJuxzWrccc9dlmjYeaGwnzBBvjKkt0r6XnVOilp0La/9LukaUG
XUhA4o1TlpzbWK6Y4g7RBPtFRcXJKc3ynubO6BU5Ye+TY8EGcEcJEWtofW8n4xwyOupbJsKJxJTY
m2czyH0/HTBYyP8O7tKdpnhoO1iWYjL05OnH3Iqz9bXrYBTzd/8Out19GkKVdwXtTUk2+FYgCnDY
+x5c8jhb3u9ezPiPBuRj4+KH8IS1ZEufK/LDnBukVGrBL6+cTyzL3kyxnq6GWWCJEZcrXIDBy+Eu
4kRq24nJ3fhT6l0lCYi9rCXpkF+T0O3Gh7St9HjlECB6yWmTEqSKgu6BWmi80+CbVaLAGtP6ds85
PfhpijI/LEClkYP2a5hZI5q1OPH2zvVHyqVdoqwQZu5gCbpVsktCZX6wZpsi2mu/mvqop+KDgGdu
3AyP6C2TIJAiZSAMS6chROExbPmNIs56YguSnJh0QZlUjGoQDBy1EpRE6UJM0pS6du/8dBbFbAx4
3Rw6P2KeaOAA2+i8Kin0BFY9JjqvIE2GC4Oh7fz9dfgk83NuVcRI7cuQ779dq4peFpDAv76biQbm
1F/oCPTCLYgX7uk6ODpJkpfWjJRc6Q69AYzfgivoQFCs1vwhZAmq0c3OFgVQ+C9Kw9Pj36AfU+Ze
1NQQHGmRjkd5uI4ds0lIdjLtDPsV3gT/s0tvZYgCgoJKtgHMywK8theyEVf2M79tulTqPkR07tud
JdFX/BbqDY0+VFOA3flyobN7QYrp4NE972G7C6tws6IC5LZaU4FmufKJaFErAl9N59fMnHlXjgR+
/lHsi63CZIc16aEFUGehzcs1mQCdLdG039rqRX5whLxP0sSsjPVb/MUYDlgRcei/kI20G6wYAIzh
gGLKiPrpF9z/BeIYYMCtWHHjNVvaP9Us1N6GJk1jlCiiaOEur1/o56vB4pJpbNoCk0xhYK3jg+bt
1XT7Ao4+Jn2dPOS+1UJRVeO/sFJa1E+L+WOKcPU7Fc7ftPHcmWB6xO6XzI7SOwiRMp/yDnFhsl96
KwO41WLRzsn6HSZ+0FXh5bA0G596MmeGp1DAJzCwRZXBaCs7BnNT1zEosOIVgddF1EsTi+OX5dgk
dF+eRXflsbojA7p3L45Ty9Z1ZY3Qnw1S+5XHdhW9iTbPyhovo/y0bt6PiC+Kk0mKDLe6E0yuey3c
ZjCbaItn0C7L14gVY8iCW9iutXeMdUgOi+go/jjfh0/fa7j0gt3hjVdFaYk7HC8lEFX1s2DGhtYv
fMFes6H3nVfSuBio2zEWSqLYV9TdJJwqEchXJRpq/CtaynIYAUdyONGYQ0j3Su8ZUaktMb8orNUM
7RezM/k0Swj+sXtV+KfMCtJRnhTvHom5xNm6/5zYzNyIQipDrSDlmGFAT1AjlIzSRPq5Vm3gK5yt
hAHeFuVETadmKrv9WnioP5kRnarv25yNhaiykh/XZIsMn77tT/exiXMm7CovjKZWZbZWvSp+KDiR
V4eYnc6cVIvIIp0CZkg0UCPH/mpTDMB5dyLMs2zyiWbf78fmGkFeDYIjdZhXb0XH71TRtCmK+x+S
dLUWrYwLza+uH5C0PC8Zj6mvBGBq6iFWuf8wRSCRshz15j9TPqkYXrSLCJMyPZ25vqcTXTT0fPgR
dshwQZne/lKpIL8nSO3dH0dBW4Z83cq77hOdOvK4yZEvOfGVy+a+ez/H9Ut+TQyNSpFG0ZsmX23h
c6e+4N8XokLNwpjI7L1NaiIOSuxO7DJTrbIbwa9FFZNYVMZlWr8S+uaLLO1Q+BzBs4O0CavH89ur
O4P1hOmJo5JglCMkO3wV1raeN3Dphlw96R44r9YSjSG8v9o4UH6BuvMHERM46+wW2n/rmXSUPRYK
yT+87bX97cx/eISSRecGNePxPVUiefVZ1oITevhWr1v+uaWfbsuAcKFs3S8KEOGo92tDm36z8UeC
Gap5w5oZHeYTfU6ZiZiZUFebs53pjk4OZzkTKkP0mIe7WYOuKp06HSgR2vvi6onXdD0NNyeSTmX6
GzxbSUjSzAZjSJrLx17URKN7koYuFFbV/wTczQpO9wR8E5Oizwvuxo8OUJi6sCOFyisVGXnbT2Qz
Y/8CG3WMMz5mwpBbPehJQX59kxC0CS5X5YXVq6E/NQxYkryqh2O0HBVgZlMsjoYnGQKQLKrUrhMm
CpRLwSYVJ3T8/VGB08rzcS6QxOG7YDUX1lxgOx5IeguqxH/wnS/ZAjmtDlnJ94mhlcBB80LLkVjF
eX5mViwiTRYa+N0HvrcWm30v0jwCoqAo53RPLotsHw8qmUraEHlgJwYquYzJX2l0jmKqqml3jJpg
tKHZUps8Zkf4BWFixU9PfSzKURgUEpEB1W17OSovRck43FD0Pw6+4xaU557x3mqkaxr7SAn8ikxI
/nhH+Pp1hrXWCz+G8AOmnbuyOAYpmqEoPrhfvB3mfXcahxuQwRAoCv7DGPXJAk2xeklM+JxzguTN
lbWWeYX9QWJkape8MowYCtjxyHAu5c8ewUbKWxnFd49Es5gzyWfPiXFuZV/ibDHDQq6mFRLdln4b
GX1QCOFdPSXIfLkhKl/U8HqjmXL5dF5UMTKDi1nEDVzgUsMpaSQz1j+bVd3Mykb17OsJCcuKDBqJ
+SqjcQDRlKhwpliHsnixPsfyjM43G543wrZK/Ry9PJX+5pdBaYEVw3wrn6ZCdXHCda98hRVw4Ov+
A/ZNi72USxiya5N/0b2oASXqnn0UqshbBa599PZCtxYy9J6WwcsoSvajRKJ4W4JDc9108DkiW0LB
Xx1OPkSgFYJ1SdPkbvTMzAHRVWIrocMqqNTCiacfKrh1BCh0+jF+tjoB/iNpL25NwOzBJ0sdhGAl
cJXt97tAajsuEHUVeteJ8kdLGGMUXqKhYnRaabccRIyS8UJKTnOF0J+DC4xXoTUsNCBVzV7cdrbt
yeH3edOeAVZqjIafpdit68ofitl7ANUupsfvkntnXEvi5ZomzkP36dQyQi9+aX5jxup+dh5UqB43
Jiz+VJCQBqU7Ej3LtFFtxtqN2Iq+ZD0cJf3s/VFxmmv61xidXX6OA9HojG5tyihpc9MEJ7557n83
ZoZRe4hNHtrgAwr14IlAq8q3Eb1hcO5byKSxT/SMPNdtXKh38t6A9OuGil0RL4Q5h0wmsp7TmpgS
3Gc2ymvTELatfBR20vrBa74gYQrL3svbi0oRhwM/ZVc0DaL5GssEAqpwjF7LzwTT0Jnl9dfhyIJe
JdejzGkOtwE3V/uIKqRBEByS6teQHR9QLn5FWLCnxyBPlwUY0gdoHVgDiEVqXxIJENOV2paM6Icw
Y+M+BKhfYvA65WmLUT6OmmdIxKdKw8B7dorqEnAJpu+azuNYbYajFRwpZXGh7S1l/pK9FLWGO6KO
y5r7JxxeJcFb4IDrRgzDB2qQRj1dAWhjT/kOmCFEuEQb6G2uOa/6CbV/CkjRa3evC909sxnH2GVO
m+t48VqYHTGp7b00u4VfKBfDudkZTUENSz52YWnHGqdEd4dljSE0wCgahKb9DydB8iWNXFuLrMbD
JwtSwagculrytV1QVBVY4WdYq7iEYBHO+qxRhuqWfvPVpP64cXAfN4k8/E89WwH1acdAciVDd5oI
OJLXIKaODCRzo7c6gh6SG54dIxCJniiB5XtCAxtb5MXeiCE8T1MzLi8z6EmkLa5Ome1tFSA1bwFT
YP/5CUbd4vcI9cRO7Ok2xfJe17xJdWhTCMdkSO+CobkUbvq1mbdOheuqNChKxAYaBvNQL0ZIt+Wa
3lRNPorhp6lmTMYmjeBN68lmicaSAbRDfL0Xs1aIAUvddr6inW8yvti9x3I+PpS94ks9P5XTtv5s
btsN968ABt3QpnC1UbWHQ7ZnC0dBDR79Vd4X+sMOrFbYYC/+d+9/QCxLxsMGbzH+KbbmymFsdX3i
GZOe8v3x/XV6hz/3/RmQ7nSBu2+MmLQ0iGAi4kB93xSBbij/D2ZCTGIF06fKivr1R26i6kNd6iPp
xNTU+LDuL2YA4QFCkaK5pjXU1vx25xcDUIUPe0fnY7NfXH2ImrzOgBpTKFwjUEN/jtv8tRTkW6VP
4ESKRGaOFLs1QT/fx1MMcekMCJ2o38SjE7W+ul46oobBcEn723PnIYV0FhcxNxcyipA6eT1V8hRm
hHZJWlhiEpLSwGqI3bowI3ESWRYMitLwlY/hCdp6lM54dRMS5SnR+EhbogQKRZpHN2MH08k5LXFk
HkYIN4KVHO+0AixHDYVK5rURl9XaK+O/STav0v3NSoj/EJOKYs0cJpSbcOKWf/NeKh3p06Es4tnR
ZC4BnAnu2xuVmv6YsdN3ayngI/Z8M0no4bHFiYX8j+RJpRG8PakvU6v6zWXNzGnJy85o15aJuQ3V
XBskbWoVeNsC3rcRtpyYDTNZ0Rzle1bUPYxjEFxA4M2nFCMblx9nRxHzponBQMPfy59lPd1vb3nm
//NWMvk7K1XFBl3/59lGYPcyVJPdDRlT9hyjAMaRQJ+wdElnDDw+4zxA7WD6+VmpGJgvEaMhGWkY
YgPAoqvkHcuQn0XumEYM02NYPtupYWjbNoJWU9pZQ0dsLiYFjwhCDsp5KY1QRLKlUl87dKChlrDY
w3e8m9+/ny3DzfJv+Q7Rk7uqyPmhD/0PENgF+32L11gyj8SLxIXZ9K0PG09OXRc2UwizFPEX9tHh
b/wxRrrwFCpJwxWfAQlHkNhFNHgcwwUqYRsyqqzZRcPVob0/1wjGNaHmB9UQSiuvYMwYwlszQXxC
Z7eZjTZsDAVZIG1SbZnGGx72lr2bM0dsrUU1azbo9CW3Le7VqHInphGiDtllX5bb2v0TUChQ2RuV
ZoLWHqa0mNoYFSQMMVZipCf4/wMmrXgpzA0IU8DGB3Hgw776DVL2GrYiP+/8IgM6i42fNCCSPUC8
cVGKdDpgQmp/g5paYUccQdEJyExQwDTO7gDHsfvaT83FdklUyvYlEnS20TFdRZJIA+LMx6u8olhf
KDJpD0zQyEu2CElpUORFx5DIAhEYXxFerGjk8ImLGa0rHeK4Joue/1IzxSolRnEAvnPHYqe3s4jY
Q2bhJ2gbRi0AJGKcyfxmRh/I2FPA+F/2jByuWgGIyGxM+nHO8kGZcshmwv6IO0mdBKUXHjfVDRRO
FnvkGvCGnCFgW9B39ZqORhrSqsfbFIj4rDR48Qppkko6Lo6p2QMp0zJ5R0IE/aJOJx/qrFlRL1Uu
sE/S6gfLOVgrrGb/RsGZr0xuGAg65btx4KtWgl1OwgCvH6GlY+FTuwHwpY0XFMNvTk+J7Jhqh7o6
D/oDddYZui8JyS7zyxS8BQLY5eA3oxmccXEKTbfqmRcmbanvm1BDXe5keFJfaKubkr7FvP8wnPC5
J9o69dlgqS+tFOq8GB58SoEzGYAO0VK9mg9awq90ehI0ckx1zTIRXS4tstC+Foh8nN4hD7qhKOi1
SUCET0ZHRDx/6Aj5NdIkuoGKxgMjnU0jTZF7Q3Iw0LcOj+bXNPDPnt2pi5JgD33ZmYmdBSGksZ9F
SWxi66a6fUTv0I9fYG9XkQZCGEWLf70lP3JwhlMr73WHUIqZwpVlSll6kgb1Sm1B0VM4cLvcDKxI
UBtqd26xkoaB7JSoWwa+6UXawdZa1GnOdbnzjvwRzop9Y6sCvEhKP4txHAz3Pldmb5Q0LKeqQ2ht
z1BYCop5vW9zfrptDgaWKlUsxDigMy+SFxtknW3DSz06jlim0OLbGwIcampuyR/3GK0FWWPH81O7
icI98gB8Slj1R7XGN7Z7jrLDSmU9fRzd0NnxGQG9C6dU3u/SK3j+lBDi+V85O0b+FL41aOGIe5UE
MXgufGS2rwMx54Qk2UHHuf4W0PPn/7Y4nzYcC9S8dv8eSAyep9XCj5c2q9ZZtQjbqfvwhK4m/nsb
wB+mScqzvMK2g+oQ+5XNWBXMT3/Wv/WY39wr+0ClY2K9pQk87yIS611F0vS4ESmUUw+ydAkMcneH
sqpGx6ViHTYNKKZ8DrVz7y0HrovWnKP5kNg9uu0fggWvGb3OeoWKgprQaeLj1iaRdYC1WP4ppX7d
WYbUulCzQjDBAu96YgaD/3++g3Wemb94DwOnfD9ySowyh47kzELwUYVMAEQt/kaaD/UcRXtpRvze
l9nbP1YtFyrpJE8UIwE+giLj3Bp/ULjy4+QF1ZdrFi5mEJae/P2dF4mzCuBd8kTiNK7I9/skSS3V
jyM3UI9nL2MRKKLei7Wi9N1QVBq+sT+MGY2zw+GPct8NBnlNoSeAkRO38nwSVtPouLdslElCXWig
01SewNkkCzgVfj8A+AyMsNzPOZMeh8GRdWNY5DmXXonPkTKAltrd5H2fLJhsJaM3e+j6WHkksUBS
f0KORMR3wiu77cL7nJs+GEPHZvzSC1DQ+/vmmnSGU12pzMjE6emjK5MV0DbhehbGarqJSCNx/5rU
HfzvwB3EKEABj0DN4MK1FUxu13tz9DcGuKJOWVc5nszCUSYgnj5mDiMuqXxDidOU2NGtVMlCo4HJ
dR2WLy61oVSpw/PGDL9Ui35fB4HbrFXSW7FZMTxrVfP1pwx5tcgNTdYYzaqghWC0yR+0e0rW7n75
pqehNPL0bemSH/k69gLsGjI75CblbqimzUWSHYNjDvpnKggNXPb27kY87zs560rT4c2znoAQtC4A
0rmlkUps0sogLIJVDTjtAwoXQ7o+nS6BnElD3RhV7mNBbPaFGyujJ/iHmJ3Zmwod60nqh3qh42Pn
JPv1lgHB9KLFcLuUbiVzaxiwqnufCHt/qUnZ4XZVMzfix8RyURPuLCfq9B0nuRTd93lEvY0U4Kgm
PSc498oUgVHz01CBVflwrQk9kKwb3Sw1xIATdtPK2uW5CT7Vrg+n+98CwVFX/5SqRsEmDGNhxVYL
IBY6VEJEFgrzQLsI4yg8bkwit9FFd1XcMjatnznZhRPRwkoXVTHnDn4CnjHebeezVp2k4sLfURl2
7Pix5rqMa1SawwKr8ZAHaKtfgxACObq6Zch7F8+imRocpNfUaxV5LQwoPTuZPdxOboWp23KksKcm
Ei6BRO/10O7eXHhepAYL0vx8GSeCpwgx4uXNSb3mL8Gd5mHa9D3cFLQm91OKVSvhU/XNmyVaj6VZ
VEVJBwGeuyWAvhrACO+QrvCMnVX/g6jqyCNlu9EGd5NZci4Tfi0kqM3pvMuEkqdt0cGOy0MI/VVq
z1PVPIkQBzDcrkuArTRNmrmNNJbK3uZLqYQg4rLODQFLNYPfhKVcRCPF6WhTufKSlHSuMXuHYsqu
aD5i7MC6BevNF0afmbqAWQMsLFEUGopnctfAx4jT6rUKSyceRQZdrEk9cEc3HN4a3hpG2zKrK/Z1
E0BhJavcvrBdLnTJUC/qRBAtl9AMx5NrXBTPHAufv0RBbkK11gTMxarQKIAgDSFazyxpWker4Q3F
wHOR5nR1gkbrIDAfGeiVeLF2EzY0dOunnOYaEKFgRoYoHzO1G195ZPjPMqGxlCXWpMTTWXkVVL4R
VW6tXKzYSyhHiF2f9fx25dbUJuP16P385+Za88XcrPENauhjC31CRU4wd7uQgIIAqjm1n48Qbh9+
epy5FVDg/RFUAbVWUmA596mLrRRMiRD0b6iRWYFUmbin+LXl7VnBpG/xXMZXpHgqs6IxT6P1+MxF
/B//T97b1Utw3ek17qRkoKDCJCuN4nub/1OV7tDdmb+sgw9qDjkwCLTAI+AFZ24Eh3RWpZs5p/89
PkQVpwA1J0l9JyAhtLSvGXKKYazS7B6Q3ZF88n6x4K8l1HGCSmnVzhwNuWgwxNlciZ4zKC48RimY
lnano+FE6vGeVBdbC1QtFybJZgdX3gSmUakT5KqxzMKUPP36AfEZ41SZ6mdSb1t8ujUA3YYKaMlH
IecYyjo6T42Gs0AZ5RlhvWMGQf3ZmZrED9GKMlPnvnc3hZZbXyYPQtHGFPIBjk65DhMY+wpR0AGN
Q5m6M/tJU2JkGEo8bLYvdO0iMpZibRzaybkj5bSDYw0dvnMeBBU0AaBzUESkxeM4QBeNk8DjkJ50
35yq7UBFU4QiQzFnhFtvqfIF6YbuwDdIqXVcScPxiBPmYiU0cp/0H6cQKR1NxQr7oXyzkQ5wAY5R
rUrtdb4wl4nzMifl/xku6dZMh0K08JiYO2jyv0qEzJoFGWLj72JJSwu3QqrClkKUkItC9WJwgVBI
a2/S7IQs3DVv091FCCVmAT6aPhtdfu9saBw/DgpqyVEXi8L52FevDlCIKqnmyQzi+Gt6gXNLe5Bj
FQYwHLSePM+5bGLxbgkW8JhNbVzgCB0uDm5d3ow2VfWeGQkaI/TM7X9i6bq/xyA7Ll8IzcoCdYzl
jYQS6NKylH1gmOpSJgaL7M2SstS+fU+D3oI/gBDqRXW0iLHqulKyDQhj1BhHTqCkal34sPw+qUOn
zny5jCJugaiM/NjwgSP/L2dXoEEqRQG/RG5b40eOxGtbgw0lt8+nJ+ob4rD1Jm6UxZC6LgCaczF8
FjcYTW/r235cAiBJqv5F0m/bSPf70BGY8wt/iyHLf5czTZM/gZNhHf3c7OW2iA2wwEL7OpPf+oGh
/2YnmHQxHZm+SViAEiziAQlPBx55YSLRtUxygN5kXpclVrRlYMeV6NXQGCz5sgBjWcveE+/KHcwx
I0cF2NTi3+im6FjKVzsox7cyn6EQU5wBCT8nrlzxnG86TLKBMGgrH10Z6dF3v0NQompDkfmm4DjZ
J3DB+srHzawwW6UaMGH1dBuiigZXyuDn3wAeFUC63oGWUOK+4k9esQoNRKSgQvP4FY92Ap3pDWQ7
ysRqQVEJ2pPzL5YihxCOh4Bjbtf+eRn6eK6aNc9kyuF8BkxR1NEyCb24ozIpjufAuO62xC1gpQ6F
OZEvWAt9GmlCeJ1ZFn5dhPGrhhjKtmA2lRrg4HgwDqaWOJNBqA7QVqqTEHJjPXXoQpNoBLBHbF/h
xCio8PLxMBSQRaQMkBPIXUbrc9+WQbd5tY1EjieTjKd17JtJ0NoOtPwwCMRwYyJyfN7Ph/90OHOF
bbxkjotKnYobrTHPZMiH+ArtbTQ41QjLq1G9odJ4XXiyZDThWe4oEdCMNnDKOhy7g/hBz6TkX1e8
oAtY7lJ6jA1bZdx1LuX/iEdug56eOgJI7/6eEu+d7KtP7BrmKg6e+y+MduHapQ476jAt3f7uH58f
ZucQ/XXKmK18FO+PUTJgPqK2raWVxjafI3Z67USeeRECtiosByOOnwB35Dun23gFFz7pqQkgSC2x
VCbcJ7OyCg5owtKV9oOFhHQMa58mkb+v5O06Qq6O/2+ZLmSySZ9x2tJ992Ab7NN0x/Ym0yZwyDte
G/TTZCtaxdFljZbGKBgWZdPSyTeRoFCexpBlabZxu2uIbNNJ78vTiFs7zSN7rOVEb94OCGym+aLG
qlyTza6YRXVHeFr8/k6hxFuFJbHtJPQyT59xcWMXPXjziU5wXDb0UvgdJFbFSa+FweHYjGoVfkVE
cw3YeLs1FgKBEmeDXiqsqXfOGsmv3yp8VkhCWjYauUDRsHc5n/XL3vWtA6L+yCg+05jaH/mI5wMT
G7SCJaM6T1EIYO8IMoI2W4Uwj7KgARWwuQ5GbXEL5pgI6PJ1bQ5NMvKs6BW9CPgDl0PT/FZtxUZs
0Qmlq9QQK3q5FSdZNMtyavAnwWkC9CUj3bw0KoLk89VW6QPYKNAgaOcViE4Mz38lHIrGilzBzEy7
uBlened5rhcOwSLFhNxrAQ1QdsAs2XAZPnMgTeejfpMd/yh349JdI+THS2wJNVCKDRUw9EQ52Hco
2b+9z6qtz29ydJOtlOzzYNLOoc8x5MBlmFMQr8yVcV1Npkf1OjP71crNsV4Mi9ZrMlT2IGFoA/1x
QxDFeGbyntBUBVC/NHewaiHMFU2gSLZa69GuNfw/KifTji/8RVHF3zuofEPtoNoFfGuHnLgVcJoO
7IjHZlEbybvy8iJrFVaaPyLwaCJKVQbtXkWk5m394ljGAH8Uz730cMKu5YIz9yCsxcsgbT1Sf2if
aUxP3Cv+iPGaqRPz9naYZAa7wSJVebVrsNAC5IPaM0MVeFLx74UDgcr6K9YJyY8d42skZA/tIDHW
KIVd6z2EcehLaArZyiuSe3Fitj2FFT5vRblGZcMqRmEos8Y9+vs4K2Y9vT0EQ6Pmg9JXI/BzNtOo
VeNOtQHNmuuH4ZqJoDAgjIXEJa83Pb5i+3FP7dBYorjFbCCeTVtsuK5mQd64kFa3RJDVKWFfTZ14
iy7KZHxuK1FNRUSeUV/u3PX0MnLBFEv8ECOy4ls5NUGpWJ+pMDDh1b9USc0LXFOB7lNHv7CrwyZu
GAHoKw15hWwAwAnPl4wVQdTZ7+XSZaCnXJadCNMT+Mkjr07+evFAd9TGPC3ELk6mbwotJVxa296F
4SD/NJBeizRKjqjmcATWuNYj3IjcM9wmTxCkFIMGg27ueYtfAqge9LD51Q/b/O0IMiDMs8AMHQnh
0q1ZzwaTMer7wkmu2oo7J0NIl4s8ewnmw3N5rOYJTo9/PR+VVS3tG3LRbaRIoPbUHtMe2HYGfjBE
A+9LNJoKBkp8ce2atwKT5NIFx/YUXaxFGWI2H2Gg54cU+jVftzs5Esm+sACUpcIM7/OqYCuGl7SN
8Fhky34J21B+HVnrdiz70vcZuEW5mGU3K+E1h6yL7bAe/YR7n0AKtrq7a44IxjEFr8uuA5REDfdW
SB65jXwA10tKAfOdrxgg2Mxhuyh6E2+zhvKpuXlqb9iV1tUGa0dohHxkxVJskcW+K7eyYPygVSI6
ZN0f9Z440/0RRWw4GVeCarOIxYKJ5eaMpsWDm9b7Ue/Pyfz6tM72NE5cY54J0zkK/AvmutCCxQw4
dqPQD0F1G9mpJ7fcG6ITSmOXK+Eg6DyRItwh+KQaa7YQKRhY0pXu3OuJrpBAtA+gOjU12Meauh5T
TnI38reVfLdQmCoEORw64bdjA6a7ezfYV5/wOvE9FzQl33+lLxtXwfzWx/W+b7KhrwxbPXu3DKrd
m87mlALy0yfEvmWryloZvla4WBZMWxkfLu1CPd6GGbVo4UI3OUJRkk8MXypEhWQM4OvBzQnQxsUI
H5gVZ2qpr/lCOeb9fdRnyztrWBpDw5OEXaHYDDRm6fzVfz8b4satgVmO0zPZyFx7u1OaOngV+F7s
321DQ1u2PzJedKIhwsGd3pIatXE1DDEFz64oHlREKQQsFugJ1wXOzR29ChkAJqCmwNb8fpnZH21s
4xe81+c/dw57u8Iv/VWN4gg6XnImyaCZ4Fc8p5Z4KdVIAf1hYSg515B5qYVEui8ibAoitAYOMlP1
OtsXqgTayrvAJmwUyCedioMN19DOXMCCu10MLqXoND0HXWSF8rhjrPLyanpZdkToux4zhH3YjHxU
OmSu9Oc/ofNCY8zgapEVeSx8WjrXa24WD8ilGX3lf3LPllk1wrmQXiK5gG1vkbMSSKEfm16MRrPy
wpkPGoaX/arGNB/kxcZ9KFToai6NU3eEkZGbH3mOId7FNIXsipTP0ToUcgf9t+3bxVm9Rf4olNoh
PyqVnyLdjtHKHKQzVx+GLxDi4w89vhri8epW2tMqOnrv8GrNRiCkro6Q74YgFRPKFQxiZCQSfSaj
0g4QwGweGslpjXSe7GbXSIZQmNL4GW1JHdevCNV+CfLEuLLfg0Wej7F66/hhuQAtMdjWyT0HLKCy
k+UvqUrKCTm9s1Q76+1rn6DCx4tM7wad4QqRKR5m3rZaMUcMOzpXg/lgBCn5YiqFB7E/GLzH17Au
8I04MWjT8n4TrtnNVAq2cfW38T+DCwUb6y2LPYKnkt5xuLlgG6BDUCT11RSVq1ihEIRxrXfyAbVj
yYDO2Mxu/7d2S3ZD90WPkucmPQRussHKFeD8R/Wiz8tvJ28dKNR70xtYy4cTdnE+yPKuyxucy00T
l/RvSz3D2T9Xi2n5v+ZmHFImYsJ4raXGYWOpMWTdLPw7BDxumWTYx074nIL39lWyHAVvGsntDhVu
Um/d8Jxjn6lSBn4Y/z58CZuKSNFQmlRTX3ZJb2n0Uytj1QNeaceYWsWTduAPv81At0ZENIEt7sHX
e1+FmOUwYfAdS3XZhevyOSoENxDrwyXNrDQ5ocEaZXL3Qmis3lDYuHhg65DVtiAH92uUVynwZrWR
63Vz9f2Ik09UtXFuqpte/RvCKSCu+IPPUIzdMAPdeZacVLoHkWWYIiNmsX5a1UsqptkScHLoyWxf
nNJ9Tjs8XjDkEFqdwrZedpEpy4ymAgQUzdIB9gTaanTAbp/AEYroqHwfnMa8BK70EBTrzVGpZvnS
R1EvYS7maP3AaqmmuW75bvWKh1mkI+gLrKpbkU0/wH/CS17YPsPWps+tTJ/9hqagvcZLwGvrFr9Y
9qLmIBbHmnn9BRbjlotTiuo5RvDO43eBk7O6V2vmeotHQLyK2rmRHZED8IYsr2EWeWUikteP3Jfx
phGgMtU0NOuf+7jY2PECJie0TrdLHCnWpfk8mqnDzxH5hOZ5mbcl9Y4lVzsR4mKPU6o7dQE0gbL7
FEGSXQyAhF8n9VbxxY+w7DQvnz2mUtiV3Pv9y0uW0MHri0s1v8XFzhFxXh4pMGjxjf3klmvPN1+P
rOZfv7LC7CLntX+nrgIYDYCvxYdQkXeDr7lkBIbA1amd1mlrWRbHooHqM/ffVv/n/4OwIIcHZ6Sm
dI1AQG84R6xYb+YVQrXhTBqFwNN3Igp1We3S0KdB0MjZry2aKaB/sZqLce6sqIVpYvrRAWLYnX7l
gjHPOpLQ6GFfcnBOQ2qned2RO8X5YK9EXEs0Rer1hzjCfjIYsQNCt4sm5Yh5lhnUDFnB4wlg82cY
bkGzMcRTHH/eqJh5S2GPWJRyNdi8d3gXtTwyhBckBjikiZhS4uZOPW7gEvUryDlvKBE8VDDW/rTj
KuPKXWYpxkYIgwhgF4s94IWOHoErKqhjKs5f7yRda3gM1bOru5Tu7YYjLda0C8Y3YCwk9BJMNDX3
kwlKN3f+3r5kVMYhKAi/u6mMZ/Ix+CdoKNCL+HhVAfZ2aviLGMPdy1WT4viWlY5Erz3xgdqFXoms
G78KzqV3KZdW3N1guGbYoy13mZR18p5fnUMCO2HsJYT7onym3JTzFjenUEpxnpiDm7w2OTncgb79
rREkKrhg1f6wrMQbAmHiixMIplPCEZ8Teyf4jb2lILjAISFIveSr/QMWjY5+Hg3+FexLzWUxhhnb
Bzi/EJ7xuAuXEC4gPgAandjfvOGjIvhAm5pULDQr9nr+HYueQvBIJIaaAm7OyQCYsQV6XXxxjaEk
XQLcJ7mN4XK+l+Lt5igFPYas3HvTk5xqRnU974MZ0C5WI9uwPdbR7WmprpY5WXJlJ5Dx7mZYFtjk
EPUEE4KfilptITVaGVf1AYan6KnsnKleev5qCXsqUe225n1l4U2N76agBWVUoSZr0v1AUxAIs1kW
7XX6mOMwFaNdzZMLvezfZiyqG5P0yDV1+/fsRPXhEyjBsjEh+LmYLpe/7wiOI1VXzeU83j04QP/C
HsP8JvCn+aXopWFTtFjFAecKtjOChTgY4ne1gs7mPy7H4Uc7Ev74ih0Ily2q9LhKvWLmOOct0Gte
Copkm+MFGiy9R8zr6wXg0j51jDwS9F/lIwndAx9g744v/j4twTORfE0GHmpaSBcvH6TzWrdXDwVQ
lyW73jWiOyEyHNBaCxuetbnMwMOCor/rndB1vCeRKmcBXyWMRcY9oqS5/YiPIyq4ukBA67qxDNjC
6fw3tDnwsTx2AIsMobMdjJYqg1LKIqVb3Wz/EmvYi3T9+eZ2DaXV6NrraXD9DclMSd+3zqYsr2o6
vkr5ylUps93NVE0rSwNMqjFvTdRYoP7f70fBeKtrrLveQY+zvgYaxpT2XDQ0PyO4KDM+5VzacszL
jU/8I6rVp2v/+XkKR73Aq6COrdr79s/L4btPg/BbtVewqiCyo/g/dbILMMsMjmc/s2uliOTQduVt
cnIzkHwCOAeEemd/jadHvGyVFYiqXMdXET2VKi6P6A7NHGuCZ8fl7g6udNeMqAvxp7XT1H+zSK+M
apQ/xgIkbpv2p9dfioPwS9+/5yNtfnz5N2KBzWpusPJYYUDeKUFRkJ1UNaW3aHu5YYkcbb2KHWq+
qPJBjJMpgNPKOM1aH3noxI4YQZe5ma6Wc/se1nslxPyNq6rO/nQxGRRVVP+XByd8IduSMLpPxV30
MnVo2H6fwEYhe5u/Kf9xW71v6o+zlOh/dUzgRtpNv1h/2XxbmhJzlAdCNyYoBxIGFVvEsDzZxQn3
E09KuoFoFrDZU7UPfRRGPP50EjkDf5zHzdpuzlNxGa88MV/CUUq5xnTtnfV0RD41H/LqQHS1Eo8w
Th60V2N5en6kgo4hrctrxZdwYHxJm4p1gtPsWFrIrfEEqfBnhA8nsVNkFJlkod+JEAWfjF+EcKgs
IfALfj6Od3qQir8pU+kQhdoksYXfqMvygxBW77QJ+EUGz1/HO588OHDIOyr2KaA18V/Q5CuybzZb
IB5c6iBMBw4Jjr5bZm/RJPd7ShwpFzUZJP03svVTJu+UF9qwNcjqIoyl+qeDC0izohgojMMJYPBN
bCrfvr9Zv9IBZYORZh7eXR6iLaHwV3qgezGKSQpwXs+PijELkYPsKOEQpytS3Zigogl30sutf7AZ
zqpLAWauwiMME/iLkuabChGtGKSXkjQ0oQuDOE7dfDzYm1Inge6VrtotFKYatq/XIBnFKidIUh29
+lkn35qoN8ku1L+Jb5Ud5KWWAjLtGKRyJlnXTuteaQCd8rtb65SJn1Y6LpKnbG4rSQNANjkTTm8e
CpaFLqk98m77Z+pKQGG3hPR9DcI7kZEQ3jd/FwQwNPMJCvPiMj8uAr/VO63IiVH+9sgONXnO6TWF
Cb8toQpBkEdBRIqml5fXmVA0l05+jMqe57pyHeMD1O4jjMurtnEQiIPkLbS0VRyIJRlF3frCo8on
ExnoJ+6N0yzK0lxNp/oJxOZHpyaqkjGz3y99xV6MwkbbZgxw60jWsxWb2OsM1HU/0LLLwWOpDyb6
BGgsfIULFJ+aZ5C+3Okjd0YeRJq6KdqVYEBHp6+wz4J2y9k0zP6KQbO9EJsYL2bTIwichjomJwGy
e2GZcAJshbAEhLscuE25RmIjOqM2oHt+2b/saKfT1e25E6sSZ7AKdG+Jk6SJ4Fa6J2hT3jYefODw
TpHgQNdt4DrC1Y7ri0l+YUf6eF9kiKHdkIMces3w2QChtSRE+MdFV8OFO215YG9SG4KszS/BEPdu
XO2N6aQoFwGpx5zl2BiuQtC/zciXivmnEJ8KDSwk6XloBdMNw1wNw9f2+q1N8IbvjZxIKqTbeQwi
/PIiJZ6Lw1IZ95s+63g7JzLcaf7Aa3TahyHDnmknHN24eQ8TQ6rxxrwd0YTVsBNvQmE0+M0/ZUfy
ZSqrEpp9FuTQusBHgyUnfmOzi2zGUCbGp6on9QbBPdO377D/adrYUetVefH+pAO+t4dH54sX++Pk
kp50wPKzJISq3VqHbavbuZPPikWIMt4M/E8fXztQPYyrdi0FmgWJNtGy0krzDy1N0hnOeYh88Nwe
IFFBIlSchcd+Z3RkYwWcUDo9SbWcUktJO+pmj/3PdMK5DTrspXSxWp6Nf7oTEV8MnV3JDsipUY/A
9sCM6tVFn5IJN/peapI3nhtBBaLKpMcrCj+KJctl8JxFbSCtkE/Lc2GThtWa3y4Kgh1QNy/n1+GE
QL3I9vcM8VunrF0SdR2YuxtdixMmR8RJoqNCo1tvgkmld0G3vwqSZJpWZ55fN30yq4RmsAiKvTgz
ma2DSo+FsY6JZWJtdzQn2/ZC5Gw1NFDl1X+4Y6d8nRUGYecJ5H/57A5W09SXsO83PgjgmeA5xcvn
JwtSBzO3UtbZZ2i4a3vnchG/ac4G9GlnV5p6d4CLh99aLwr+zx3vWZ9Tw901uHJ06Kd3iKgt/iYD
Yh7g15TR9u2wEeJI5+2pqHcScnmzSsTfeKwzuR8MXFvsuElOmtJ4W10ORkm4WEBNDTHI4RwRblIv
5N8pSMp9f2M6t/GhVx+jSAo77xUhfa7l07v5N3Wi+bsjzLgzHACVsim6wdEuSVGcbUMrx1Lo6GZb
nF0kC0NkrUDMt72RGO3vn/iqcuERmqr0aDJe/z2Ugb0kHXp9cH8UHaS19X/mcwE6g8HvpakX6RE+
pyYCpRtFw/DVJZe2bkS4f6LWxhjD2O6Tkfh/W/+JcVAB6avpbXSELup+BCEZf2q2x255ag0T4QDm
nlKQUXT0VPt/vkaZlvRuJZaocKhgiCRvCYfdzQYYUX9QrgIb8pLkEwJNHbAa6vAopabtq1Uvgj86
NDwpAbb8aJImf19oBqS/9jvC2j1cmPpfZUNK/wOefqfmlHLqsmPa0w745Ry5OGX/jn6ZBDYN8aF3
9f9t4jnb9BqmP9Wv0t+q8r5kLBlaAkjmLWh3htXAUHUzUhHhljnvo50nqNotTuxP9KH9/vC9thwT
/SBSjyte1lh5t2GmkioaNKccab1zQcL5VGZFeuCugt1Qh42oyw0zdlFnj516u7f0EsHXz0wHadZP
qU5hO76AIPXevlaPqgNN0aXlOIg43HMFvM3lPTSioQe6SDu+GtG49LvvIkdmw7h11mIK4K+qKql3
Pzu+Leisamua6HYHQ8r9Bzuu4ZW4dYWluQCrCM6ufRlsV6Ul1iXrhtmp1hMsR3CfQRahdQW4qr3J
Ia9U0i1gLSXZQjrCKBcpNvPfd07OB00XAtTth8UWjFzJHmNrfp1RTrPvobn/NP0gEw8zvwA4nwSV
2M9gcb9AMCbYwI0UG2rRM662EJoRHnQhO3RVwvqHOJPpTkqW+oKtTDNCaWvebmB8vh6q1wxwqA1l
gyNfigD8Dft3adVP862rUoZ7Hpy60r58IsvstnVzg3Qz7U1J+nBFVuCVY1QVpmpitSyAkpi8ROnv
pilWHsIgMn2rI3Co5HPqS4Vu718eP9hkp9sti6olYh5JUfQPObAn9GodRaqRl7LyqlTjPqzLXFgu
Y6UraDxHv+KyCokavGIvTjfMoF8s9rx2ef+cN41ELSMg1nuddK8YNDEHTM5LhaFrNVrqOhTYNCmi
uBvJitOyS5zVLkjVbrAKHiMnh0d/UrKc0rxWG24nnEyTQnJJm8J8vXYH68S2Od9AeSReZPXHgGjn
JkIln0srL9pSs8XPwN6P7Tb/pp28gSLe8Xb8kUiMyuMbQzH/URZsTebzl+R7SS4NbdgCUZpAKgTU
0mMcKYGXp9PIuuXuEv1PLNFOC4+aZwSkFPe+TP43nskgrvyTSgGqAIVma3b5IwHvEB3SPI6cj//G
ZN3yKNoiyYyLsC/Cssk5c6CaKBr6UD4ivV6K/PaU06dkKTlD6z7kxy+9YpT54LwL/i+JatrZb9VT
Vc5r6eSzQBUjNWOQ8ZxR2gYQzy9/1A/YP5eICeaXBy8tD/tM6+xJdYFDX++5bawQi2mOakNh/e4a
K0JjpJiXfsBpaypt/Eo6HJOqQltThcL9Ak2/6CFEjhxku30s5q6/x4d+BWRKmk07xnRSckFLHzUQ
1wdYdBOsWNMilIyyPYXaKand+htb7OV3VlyYxKGVdYDa6GnLObiM5onYqxS5Esgxlxtm/BAID8mg
h7BS2FCD1TQuw2GVSLs5LecP9usunssJHHYMoaNuAzr6O6hukvWjpFADtdlAgGuKV/sDdjfdQlZd
XxKExt4Wn/YyyWO107Vh3YQWzH4GRu3GqW8ayuLqZrMrzoGMchk0xUnPRcvYXGVYlaZ/pycpLxES
MQ79gThMsNfrD4caUbBSST61g8jovJwRA4laLC3klm8X21THM6LL+LsvlQo/dfRgLdEN0+F42vWX
VlGK29EL3KkJZUq7lPg9Aw8xR7TFV4ZMQgySr1xTwmmcuSMr0zUyK5txNvyI3iwTjrpaKRWt8ohE
KGty1hMZC2ESX7oQE9WpDndJrlmOZkJiqoXT31aGQDwOwhJJ/wpaNhIZooIqEj00LA7f1J9AehTw
V5hKpfjO3s++apao8tUMEphvzavqWRio9BZBOnRHKjgsnNE3rwgEGxglXaQkLTnqjcwAraIPAHOD
x/vRya2Y21LFHaegSLEyCs1sisZGsBCVIgRnrhbtbZYjHDzWYT/3Qse/gHACyXGrqg7+R9ow6Pdn
vv+TapnhXmKCKkGuwUKc5p5V9B3IQJ9XMwUJcckSlp6yfnN1bzzUh0xNt/2mfxhE4A07nrECny7Q
6mXN7WEmshahLcYl53stp4wpU2hrctnqH8Klc5y3in+WBL9x0WW6sdn+lKjpYquIPvgmJkh9sQYA
hTTtCzTrOf/w+CjiOfCOXOG2R58KJc6GhlmsfvY2DGBiqByOQHLqkZ1AwdrzFcxDUv2QSTZURU5G
R2dE5epW5ZEubaGc/KyFe5T7IwR32/I95iOf/COXZCw4sycodnKJf/0CBFMFgkG9o/n5uzx9FIUr
F3BmFi4nEC/cVMe975GcvjZBOxNixTIjGmQJdUkLCvUKkt75YoZcNSW1aZI19HYiPVOBaTqcQOvf
0bgVNKI20RwqlWIewcwq7mhctOA2gMi2rPwQcCw5iRdbo7NV3yRpo/ahRierun98frxSr5XBlXg4
JgwFiSNBpSGzpglh2xHGPemCJABaEXJ+KOzDpMGmGWDmkj9NKZln/HsDeWZiElte9gOkKt7rwZ+i
/Vzj4B+IBI+u/A5glphuf1EszP/OZYIo2+KNK3uixMehgwAjNyXeMvFEXlDjc0PuSlDWyHPjlLqF
WSnXiZ9UBRSYyHebcmnNLObV/3wnlvcgrLEJ3asQ/yiorspBz7DwDjIO8860uzaz0/hPFX4e5rob
bhhAGESzCuPCyoQCIOBKhxLyKjirM3O1mVKkKfpVxlLJlxWgdk2ktMbJUmTIrAOLMERfeA3jKHWK
7+Pf7IRvq5/FCtKlS9oWp4lmHxaGlyO8mqeU+rBvbMXEmRZrYOoymLl63BMWyjgw3+h53KrBZwYD
0PIRZ0jjFn92hbQMC61q9AmTIFbzKM+aZXWlIUoWu+YQqxYUgeF4ZQCIx7MIqN0GwbGsN5sl9wtz
AdoOCbSFCwjHomLBeC+NSGJ7cQHJW1jrlfOS058cb4JElV0+XO6uR15FcfkfMFEsjtdwilaA8TdS
v5QfIE8QSv/RLI5N9AlpZ0PAUxgZZA1IotiYW+EHrmCMEhdHXbaaitzPhmiMcob7HVC3L9XAEuIm
gEx8+M3MGBN+kIpiXcK+nbhbp0f04kSpzudpyjGM8gis6PIPFQ0YPB5SV/XIzpVIWEPc14+BjFzY
nc4jejZL2lva9dJXHnmHHyIXzab/SY0oGLAYc0xriSe57BhiV1CPvDSsW/BwQjxVTYWG1nsrR8aT
QdEODD+dl2NIFXBbq/gB8JEBfN0CfHLETtjjf6K9lqi+dgeB9O/spNerHSHCq+jmxFJg1hrLJJxj
sn8EwFxC8tgsulouZ+XxNDSTiGNfNrKhHpV4uTKTadBg/eUL4heKapNdWBVvU8u6CBSU2zEHLgwO
SWe852P2vqb2RAJPw+mhayaoFYbFb6NwPA3dce0uJwZ4pQeGi55QI2Mo7zLoWFk39ocTAI3JUoLl
1PUa15AD9SDngkq71PElO6MrGbndUOtra1NqSEl5ke12PYHFKhzZxvLXJ9tLRdn0/T0vxEy1VWF6
ztZrVkeuZ85kOU9+yhe4ZojVeaWITp8dSoIi6m9EXhC+OnAM1Vl53vveWej4rh9hGHDrfdgzRvK6
m6RYB8V0+jF/YwIlpy6rvs7cYqK3AGr6Eq75BP8GaaWWTP/bLdKDxxX2OZigMfZ+b7XHoYdV9NIK
IcwyWUKoawlKPj6kfAUeXMZ1MrncSvM2O6UtN7UUe/inRiSMkK3Ew0J7BA0JqixkW6yBDAT+Jinu
87DiMz0KjwaOBHIu0iIW02eslDm9EfllklHUGsxbSQ/BpTNK5SRUjcTwwyvOyEi31iL02iCvFJhw
gwt8rBbqX8b8ioUhSnZ4x1Ozm59RRqWeBpx1HgXQ4ARw0KpM3nddxSZfGPsEtLxJPZycbeK9NiRR
BA6jyNHQPs8TJ/a683oXoiPK/mZAeVM8xSQL8GmK/utnMWF6ZTryPvHvBJS7BOOP4tolFIK/Yhgs
U1Pgs8wD/V6y9fY294L2yJHcrIz8fcO6SJdGS7NoN1bvuT7GuVe3hArrUWTO3WiVwZh9Kxocp3Ns
e6JNBJ3LU5JJQhMQCHQpM5CFrJ4zHHYnKhlHuXxsdUe0QKEyfdKdyKiI/kidxmpb/0R1yz3xk0+/
UySLw9vlAH1o7GBjlyO6uYINarElTaSILEYJ3mTu0G6IdGgJTDcUE3h4OxUJKoBziOojQgvYFo9e
/O5dbxiE/mbFbMtWnVaOSCa1Is/BrfT9itECB7DmlQiVInoedDeWfLAuuBEPQAx1ByHnVnVuOqYn
kUui4ZgY371/ribX31BqpCfUKJEESdhAuQdsQwHuOiz9a5x8i82aAv+R/QiDU7lMdh7q5FdlVX3F
ieNFXsNO6UlXRfB9reXhaQM+4sokSJIWQ+AVc8JzQeRfHKb2FCqYa6EQClLGxt8odHwbzSyjNHGm
i/ij1QSrY1mbuFbx6e6JOHn9PPtXpcLDFzVlCj6ztqjg5n0eDZu4bpWOo7hIXhxUlovPxKOgXkCS
qy67FfYHCcwmmfrPycZ455wwIf+dh3jq/mCZQzws08H1qPhniXzlQy0Zp8JLYcxliJz4xr0qF+Yi
OOSoawnlGxUIlCw4YUu4Y1koo0E8zFhtpom2PrM1xmcuSXdAusXXyFC31l3uJFlrw3hw451I3HLS
vTqKLQvr627A6y/SneLJlZQka36zlJFEHKhmckMaQz0Bkxt6wQ6SBf1CKZBW9+W6EmPi/SO77oEZ
vyJHc+xyrrVlYcRFtusQRThqdXhNt6oujkviiN1BTvg8hwdLHChJ57WMrx1pvwlvyWae7LyS2LS2
lsAlc69K0XRpOVPF0Wkmtn9piuUsjs01fF560QFaliaPC36Zs7tqyy7nXhPK4BNbq5brgmFKv0Be
NHzSJrF3OerFena8TlQVC2muuyg4oj2z/kcO6DpDHjgCyBRmN3B9wIpMe8jtdZf5jOgc6ZfjXuyx
Bkrlhi4ROWmPJy/SHy0iH/jBfFh0+VyqRXiVWrMTLssruZQ54woPHg8y5tyC3S3IK31xyTuxn/NG
p3GRl6VTlRcsuHLD4xB1hoBerx4Gf0R5JWQ025O4Xuked+iTcZXik3w9Y60Edewe38zlJR6AZ0ua
93T8X/dfVHE62EUJNJ9TQcWCHYMffdV07CsMay/7aYpxl/rrqrPdYDWubLrQIk2543GmxT6eQ2US
KeqHjXpLshFrnASvzWQ1lVKhBOZNWkBrs6tvbNjlDOH8nBG7+VHlgVZdAM3HU2Z38QxnnJmU8/zf
UKWFBZAwFeJEW2WfhDUZzlP9j93lz0Zy+Pd+oJtrALwlpfFU5wbwFuVSLP7JeW8lmXpl5ej4Qu+d
MDpafgULgjZ8PWEw8WvUacdRaqD7cbOjbOnk7T1djDvSZYlx5wKg1x1mIQlJddwdzoMgejtcA+ve
C/2hPee9wT3qVIKscfy2Xk05FN++0rCPJtzz3t07pebHXCIqfIn8Op4zoxrf0R+6TQlggZNiS6TM
Aztzin/DGJ2Gw3s2iywcNtA+7WNEBcoBnyVY5BgCLwU9gK+reZmg5kqLpxrWFAlEwN80+IU9IWQp
f8GK0SIoP6dpZSnS3amlIdRollrT/JBSmqksSpFC15CdZFnL5idnG7D/GigqWFfp79qCDdBwGAgs
hoHWAXfkCE4CF/Cbdu0a3gdtijyxeyhQQL+QQ2no5LucO2IxfPxEktgwLlFQJm8oLeUtJDnqpPma
TOzkHjjpmGtsXPzCu4Pg9ke2aD+0SHleiF18dHRpe1XZFiWr8aPq7unZlCbhOf2KsaODQiUtZha7
jIn3UMSpxmo1HzLO+wyx1Z1nxG9H6oGW/1yoAHPUuUndwobjCUjT/+oKvaVDyHd6BBH5pofbHdcf
IPz1QRhC79h7/5VnIdOzpanVrtOb1cbO8fwwwM8OD49fRZp0trSdxKMmzKH3EPg9zhfQHh8Ho4Zr
aTGneXPhfmj0sQIWsIGxAHchxnw8xYCy6ccGijuN1y8oz5XyJ8BVWRK45AvYvH/3kX4qtBv31S96
K1LaF1SnI7dmy7nG7kDt+LM+oP9ITPmBIIDJ7Iky/OG13bpdnoksoD82wRPGu6Ldfl54pXnLz+9z
cyRFp/aG4x3TeebomatKmnbjUCYBQMdqJA2q9H6ECWz+uLpBfcax+HeO9ZwrG0za1JZsspouGsm7
bxIWA1bsT+Dni0KOiXrX+NVUOaTCkQs5y86NeFSd2OxiPso0uYzWP8CJQNjszqA2kFMKNiKbuNR7
YwLYVaIkHF0FH+dAdxRPIWdW7TQAVr4tgqwiqcJWWsN7L98iRlxIeGA29bqcRI9nltaIoqBjciJu
I6UfbGWRy8SMhcarvJHPNSoTiF/ZcD1EVBy8pl9eW1aKr+X9mN471ogRByCOn4PjAyWUTEkYreFv
XU5MoFt1HGh1Eyv69PoIwadxqHVwkkYK9zU0IX/dyqtkKn9BU/Q9C23/8M9YXR7Qg90DujkIUAjp
CFEuk3h58Wvg/DUQe2RL+FDbyt9kRbsjlnNCarXiNg0fRTmtc/0fEV4HzPxIktL5TLe34uEGmC9Y
u/uGCoT+SsgFabelXhwscMSDqkZjsmUF9KDRFu666PbTWqv7bxtwntfP4ZIC+ehFuQzFgGeJaXma
xJu3EVdrMnEz7Vpx4TLGpnaG/qYmRlY7BWfdExwesnd+YnUSVW+dWIE7OEiOmLWwghlFWb8uPVfK
cEH9ltuRWABEIiOTRTZSsU+VL8m3grq8f1NAatSRuWF6V52dVUAq11iPUUi1rB6kxQBSGmqesnCD
9k4g6M8FTRnoboYGlwCrJwkHX4+SIBi3rV8FRccz/fmVAuyciHLLPR+YVOwE9IfO7SqbsYS4eOUJ
Dwjr1qBRHT/ncrigulFB0YNdwL6Wj9Hl+UhwvkdYlO5hRbQ+9F+V+jpvBqbZjiGa0qvjRZq8Y8Fp
XYaohFaGU7gX3G9X7sqC0XCSc085ACBOFQPDEwEcyfp7infhhwZz73m3F6I6WYfheQ72Q3WyY8ZV
2N/aH2oNqTgyamoxW9785qYkFnTOBJUnsz/7MFnmD4HCcEUxqv08AyFA1K22jPrmGK7Tyzai+Xjy
vtLBr2NJxUUnT0HNVa/Uc/JOyyZo9FCLJlYjyTQJiIRUTlpSNoYlGCjr9hRSv291VPdLDhWsTGVq
HjtAIJcBTy32tuBaWLkCkk+CJge7vD3a69VsZjntoe9yMNSfui7c2JYMCVx1AGGcWezlG+73vyGZ
VTwbne28EJizjlfRtw3Mwj0b1uNmbsVPyYAKCXm/JuAdFyY3Hnh2pWLvhdS33cvrCiMFXmtcawqy
lof/XWJe2civ5RpxhXdgqJ4X/Mv4HH1RyABwYvvv11Axu+kXZy3j+a6N7r/w8jLVo82r3dM7itbI
mHdyl63Ztv3441yDaeB30dIiKZBcu6R97TYMFBnwAXRoy/gEHodYq8i9yc7oxQMUpth9qfQ8fV9D
1KeQUqn2j07RI8SpQmVmnhlqlVMUF8s2U55tco7ajiFP5f+cQwdfnv2821JOZoqo4rV8LnOSGVXX
tqGgfkfeznUUDo5gPG0RruuTwjePdJOgC2NcQktg94mpXQiDdx4EmttQKBsu3Wl9a5pA9hW8x+/r
xAjKBvij/U/2AFnK1TxnfI51rqyhie7st7/Kjz8JUM1BRInI1TokxsTxDRHjjBqEw6lwtPBvsOUk
dWS+DacUI02uoLvCzPf7tqxBy6EUEgD1+oAhDT2Bjl51bjXo2s6xeofdWf67JcXtSNqmQwkA18BU
Yrd55MkAsE3BzO7mXlKB1ZXq52ylNLvrGN2in9H3Vrpal2sRKuYsd5oesao9TrTrEcRJyei7KMnp
sTkK2+h9+Yp6tFfKJ1+evr1csAdcnJ86iAtNCLEFm/q9jwecBnEfGEWRZo7194gvFQyhxm0Fm9ij
5DZ9ibDijY3bjaVngwlEiY90CAlgnuP71Tcpy7ffu55ymxPz0MX6CFcVdYfrNzynn7LHaZ/V/pWS
ynRq0I42Ddp2iFrx8ToAMpaNHXSWKkABhRSmVqghT6TvWIaIKvaOYo7fyhDImQFiLu1UDDLXlCXX
ddUJln1ZmVfEo67iOjGYcibZ9A3pjDVMgRnRpno1dIntHWs4ujxPgn/OLDpYRFvba3UiPFMLAVxV
Plxri66TxQ2ybr+TVWxK9tfO7SLut5hXRpY1j7pbJ2mGjrp8xDnwwr3Cp2S9VH9dmalywGJ+ote1
1Hq8KRlfKPjbM+oxuODryBnCzT7GJLV5Xn+ngY3q1A9CphryhgdQPFuUbguLwRYc7jK9Y//3YtzS
h6JbrWLpuUHgwCuZR+kWQjE4XJzkUNrECTrZFm0gnza+fPFV4Pxf2TZq5VPS+9gWOpJSkO+/5Kd6
xpZ1ABdJcfXVXFSRa2C8KiYAKrsacgetNuIubxYqn06BaxxGvpDl/3mrxdo85WV/KKfq0lulaiNB
X2HueEC0gjVpSrsgE14LwsCWaVdOvIF7/MrftYtF+Ly3rRjwbOkt/pUYi9G7lzSzNRWh64T0aTWv
qhacn1QdY3QPLLuoHbHU8t7g9MpDV++gLUI26jJKuTIGM6ZiEbBH8EwK/10p1Ncbho8ZY9TC+5s6
LusCHW3NIwz2hs1bhsPLFp4x0ZwRHXcCncTNRUYivLMSjYU4K2QBIlqrPVc/7odFjHiscM7GYnKF
hk/oZKorVOO4rq8LV5DwWrp06d/zJ/5sS/8YdYZ1vZZuatme9lr8P7dT/EqGXRb0sIOUVT9JRVEg
7JmQ/neGVckMcEJ/X3pN3danjuXlTtlQDuI6fgcSTZwEeqhE1mzb3NsHBSr06iUGT3pDEyzMlpMH
t7iqt6AAAvf6c/9bSNS57lPJ3vG9E4eLYXeNfIZ/GRWSIXy2iEz+FNltAkXHLhyzFLsQKEsiiWiB
MzBgOceIV9SxNj5OSe++z6RAskyT4WHmVTJA4/Ox3DKFiRboLKP+k0yMnovG6rHK0Bw6w5RqLH9A
HjDW2ECP025KpkLzSYtAsfdUthbjJJKWI0cVXIwub6MbWtxAu9HX75ZGsSmfWyXqu+56H+fuLoJ1
MPTMNGKdwcmO0unubCsepcHTUlXQZK/b9JyM+c3syeCiXLuv1hpUifRCA/Km7SjgYGrTCgZ9m8LS
rsooy+U8tzmy5KdyysUTk0kBnn2mDcw+Ne0eGFjNbxWPnrR/TXpgMfyUAGih+2mfoJNCpP/NiGF6
TRkD4zi3GIu15t0fsnduyV6HpHAdc8wvqz+D6X7Iu2219ZEGLjac7neDtCVdGs/ssEDHMarrTiaF
WCErspSQ/tO5bER6lXUmAV8kL92mXSQ9sV6PZQ+1sncfCH1da73c/ilXxEsE1Qigk3pZvmM74iGD
U+cyW3zkHocrdbEvTJOrjIYoo5Y18MhDon5UPvz07I7zQjdxweBSW5U2+wEBLw2TJh28Px48soun
PlW0M0nPc8seZ9h03RdywOSCBlHmLjTGbIlq3zE+kSCU9dc0zHlJLeGANpa9I7KuqN7uJipu1s13
EZSMrrH+G9PVk5XRalUwZ7Cly+ZwXJThOYJLJDntPwvZTr8PV7MipRidXIL5fcFaPaKiCcMLJeBe
74EhEuhX0pxRKGTi5PAurMWgD44W9iuq4ENAGB2uOSPsm4B11obsk9DSO1WO1tBmMf0ccEitPhE+
igPTuIdj5B4hAHWUxPRE66zaYAa9XgOKvni/5dOQYAzrzqSMG30z3JsJWPryUEgjYcbJbQTsCg/9
CFLjr6tZxgHGoVVkxq4lrZ3612He984EUItCGOeLnJ5mHd98EsU6pNqSPO0bdiG+cT231bRDF6Tk
Y6QEpLLkH3DfokoYV7MgqcJ/UHMhB6YMh7FWtnITLNTxjLhzLkN6FFEaQ8kP58r56M+gHEJdQJ8r
rUsd5BzGDrE1uMUAs8mjqoCCEWHp96Ydp5pfKy5LLpIqw0eR7MSZKK9FnBGNlksM1Ho7yf67yPry
89GJxJQxdPo4FQ684cdPs0Fe61p72IjXpJHDwz7ZOpzXuv93FuPLU+akdBBPjNtVYFd24BnaYLzi
9m1oRPdZXX2HSXTxp7d5Jx9G1Xl1aVQuqcyIuaQI8J/xpU5nDTFGJWbLlvOIrUNHarxvuYZcbgrg
2X1xJomJIHJyEoWKMnMgShvjcbxpe1B260UhFNOXl03RLrfq/oMmCsDZyM2uM4rF51DektI9HUiX
qrUNITNzfSCqpG8jcx8Xn5/MUDlOFqv7cYMEq3XLhXm5OAxFRkAsu1Z7G7VjPdW/0txgU+NRh/Ff
ku5AZ79XPQD7ah3tOBGxzxIjZ/7cJQdrttNmsl9YDDKsEBPCiQ4Y6TKeCGqNpn17NWbcP8FIu2HX
enN+cydwkN5ElRDqOEjnCHlkZDWyZ0NXXP5d9lxJQWdgp7kAG2WKeWqxbqyB0ApIvTP0JDydRulK
9KYcbeAmdgqIuRqahe4Ro6ibrBmn1Sxd0mJ+j/UCzms5nyI79OZarAXhKnTkmosx5/sLc/IDhDaS
ZqAZ88DrxYkbK5wdB8TbzB+iEfi457xvOSLStsOArtnifg9UNb2Ecq53jefzdPAmAJeuEA2PqnTl
z2HILfGV2iHg11w+ekN79jsRTSetFn+sjrblBNt8ZHwe+I9YoS416FZlYw+C6RIAi2MRc3DPLkd1
eqPZ1oUzzdERBT13jHqRVp+ZSCuElxbVQfxBF7O6bkiRpA7dWk/IQeUKDk9pq9T1m+/g7NwxwCUL
9/WdKCeLV3r8K1IdnktoirJpvWn0Dn1bMqh7KMQ/W/ZzSejIVkWAEOuCzoNHUTPl6zSg74pQGTo9
i9KGyuN6As4KxjEQvQtJIRY1xMXTxwpDgjyhRAx4jlGZQxn5xip3w1VR4hkn78hEm8J0/J5mhHpC
9CgpPlot1bycrczRRG514iFM2ly30n4VF5XpmBOcA3xVJ8/dUx9McwD/iCPVxwYtYaptnAlCNwV4
Lp/hCDchfPXDtuSPKkhnFkXmvO0kTsUp0Pd/FrGT4AwVTBOFcUQpReVgSv0D8GKf6DPOdDzzbVpU
EdujiO3IClMCJRC+1ILcaVHsnugJ3d63OXnZ/kdGnOOxlUBdrY8hVKFSaIWt/a6+KlAZG9RRahEk
zmeXWlmzhlo2yfdpx6kHgKk+0cTHYpD0kPu+ib0lsvacVoNAwkZogu5rghBbuEBFgimN/nUDY4oU
WGCcdyVnW/b9cfwtwzBvWK2t696LdxP4/uZbA5G+HIe9ETjGwGqrfhxek4sP1oJABggcnfzFQGd4
XMLElopNwN+/ezVwblqFApbVduG8J0G0s5cpxamh83jfkFUNJx31Wm8xCzcsLUVpB0o4bADXstaD
lB07OMYqX02pWIxW4dmix1htJz+6sDjQQ/ud6FMFckf5EJshi1Scn7/soPZwxEiJS0JSQt2mYKXa
cLh9elsFFCpqb/APFHAXOi04pV8jc2hoLFZ83YgFg6B/PKVJlFBN5mWWiJwOhslBS7BY4MevRHpj
5GIJa30KK389un1crTqK7FNtij4C9RMFr/QZJpdzlaKpc2AmXSrxNvYid140ZHTTiQ7gduubcWmi
+7POgW/dmmOwb4oVpJvqnIHs9v3henJv7a4zJ6mvT/darz7bW/zV9CnI//xzQ5dl/Gc+BSeG6vta
0rNo7rBx6aBmjehuzSrICwga7/b1EjXLElTlzc/jdyjCnaV4W9nBm0eAGncv5pdTm2xHTpTDG6qk
vO03opT5iaOgM7GtOANEEqoSoTN4vM6nT6yt/vZC5IoTqVuvjUWVOxMfk4dKG+hObfvkB+0F2Ggm
lYxBsw1atafOaVeV6i1Wu8LqQpOvLF/fTqFezqgFVaryjmpj9XORThp/gPjRVNRbBU5faoQC8aAp
pgBeFztVyiocyQmKFp7URP1q06BVj2K8tTB9r5VjbZf6Z7CvGVA8IUOXN9Alv5vkXRMpxXuHZBq+
OTLkspKrJspdY0whOqPWy1T0mTfz+ne8UGWmTd0yFp6yO0Xm+9zf73YJ60XJOqplXAhiSdN1Pcmi
FsnWmUqQkYRQTBCuKJz1iP8WDK78hMSFoC5YBgXy/jE295QqDydwPLZn6EdbQU/+w70mKuFxzy6d
RErengXiSfHVlSThNu1m7x2UK55yEAtp4VnLREQI2RGSkKlDbjae+KzvXPLWAfllplBPty9DOA8f
AgfZOXhmeTedzXPVByYbw+5AFx92oqsPFFaf/Nv5vuHM3rVFDAtKU3E5a17XanJLIxWLX/gwW04B
VJfzVftKNE4f6Rr28h3ce3dTep9wewY4ApTWnTv7e8JUi86Np3ZTGTCS14OP3ZCfzisjOmNGOnXE
69Di1sDLIhIPqh4lKTE8LKUOCddOOP299p6oOPJ61ifcU00fqlP+5FTgAgH9ieV/f7/W8RMWULeA
FjfEcmp32MRWD1WNUgliZVbLAdFO7dY1z4xiKPulsnRprfHgqdIoaSxAsJKMq3hj6XAQfJPDBd3o
os4xMYty6Vr1myuSVi7QBDxDMpXRnSlCiMaCdhlGWU0dk+sHBPHyQSkkeMpmI99kHuDOv8IVTVqa
zbifbjNAmw7ueHH8vmnqp7/LeveDba6ufBfKkb6BD7SwZuTvffvwIJqrYCgXCMjtE+OANoRl5Iwu
ha1M/VDe0x1IByzXXR3BUY3jnSLFKOq57ZzwKr/SzkbnrINFWKIr2LudTxoiv+9Z13lrAM+7uwry
0W7QObx2nIo4y0d7HmmEiXb0wJKp2JS8rd1xISlEqIVg4Rs9Ivbxli6Gq3B3Fh2ea5zim252vCXh
ShPiv2GQSWXj6W03nDEkXJT/Kerxb1BlnJcFSlUwgT0uAaF0yehD0m2Ldk8RKTukYHVpDk3Mf9nb
KLSM6ynXVekE8b5U6i1zWVnmZn/bb8nOv1WTuqiK7bbDYNIOgNFvxyrtVznNeA+NVj1TL1S0/vZk
aNUhi1uC4wnlWNmIfie05pGvgezOscUX7lRrNI1J0+nOrQj94TMQUTnEQL2NnvE/UJ7AoPzUmEse
KxD59duuMIEuM3dVLY2XG3oHGHy5zl3lWdZ6cd4jdzBxk/GWYOGdtwZfuVdzOvqdOU8fgo9G1paO
2rKl5A64ALeChOqWnxBP5pPKp4DwOF91RAL3yn4c+K3iuPkIT+bvxF4pnRNmH+7bPEbtQc1Z1k6/
MblOQgkuII/VS7w39kqHRuA1WOFtKdM85f3/YODbNgeEiHK5qzL3OcrczIrThObJPAtsCkrD12C1
3gAms0plJtEKvAn+lfMclYbcdn7iMbmz8762FykiPEpmIa3mRTbSZJB6D0ZZm/FGcI29IVMolC3w
BLjtq5wFxR1+jogxoJRzsqJIqwRloQKjSBcIc+PjuPy47IUIWPp4diObQsH+yGOFMdTMuYFzaHMT
0X36lAyRIrsJu4meFuPCVU7uUCsXAeqEyUuPq+dw1RDHtfg/iIvViltchhU+0LR/SPmmIWfjq7/9
Ls81woe8XBN8370IbagvdWvXTcwa5vuqVfyTsz5QhW85KoyvjFYxitKe7tDnEyqx0vcXW4+8638S
/ulrLKIKkwUzoA/q6xZuSl6aYuwr4Qbv2xPW5EoEMPh6ffcs/nouF68MwEGAZnBI3Z57DLQ/m4EE
lqTjd/NRaVm/sfHDso0Z3hXh8TAkFryZLrLx/ZD54gqCC/gRKM0DB2vZeWuycApx7WtNqqJJW27f
j6SWxWqlb+Jhs2JY1MH0HS50b1MiaW5UVo7l1mowroEUQo6eWsfenVMlf6RBjqK/05w+BB+gSpVX
HHeLT1pfahePQY+lW8HLYMdyXOLhsu9KE6Zbk03B2sV0viBT1Yk3OhuuY8PWBQs5vIRkSBqyfHWB
ObuWlWqYIQ5hzD8DTRpO7Q1ZlsU0R5jhoLwh69gpBxYJECfWPcx17RgcOSrOUeUwHcTs6VeU+9Yg
Wy0M9x2A1+4H9fUMDN8vTDs3Sh6FGCCW4vZvDwQh1luo/NUs4Ubj3/MpdE6dQNXsbGpNcDLk0kSR
awAE2RtFL1X3p60fJ3spVA534fgCJ5WaUbBpioE4HMZdQXJJ4hmeyFotGODKSbEGy6uqnuS23Fed
gGYn61kaRE0QuxLLLX9LkxjJGh8Uzvz6eta1g0JDhPYgrzDSNeaqCV547gSA/VuULyte9/5TXqmX
iGxW6YbG5zefvpmTHpRY5BQZbQ6YjwfGATvFKecvZnt5bgyQpWUgUTNUCp3gOd3u9TxnZ6aeQ9nY
xvYLE45hooBXnJ70zMSMoPu7YgGF0hUErOmDUxbayfilf9S6vMQDTXTMuc/aoJYpYixQKUg+NjbE
Kx4jD72EIyt9rnDtSxVFvQhlfY8ynmKsQRPJTywLoHQedZBf5zEBYqe5/Tf+E3gi/6/i+EpRPXnY
OOYrf+AVrpvZp0nlXoVFxbEiYW7yisPRrUaszo9FmR24i/fB0xPsEdypnCG16ntSpu8erPCanmE0
kK66DaAb5Vj8YXsVPEnLe83+9R3YGXCEYrONraajm7Zo7D1vFvOUaX6CqeORHIioZkAk6gN+IKmb
9L09c2ou62Z53rawEHm2L/i83KZ6KJSCEQ/AWgoLYNh8geB+QQ9GLQOK9SeEpjBTBmrWdVjSBRzq
XDct3bQu3NOHBOPYR95VZ7fS6AZzQU4aYV0vPuLd+66boz3cFfiI7IqNQl9xFP7XHnaZGvRFJ1/l
8NfPFOMc8nGDIO8kY4C7eJpU7EeSIaJvL+aFNj5F0k/ODVjLyp86GI59yWUABvz4dhTcX/h1DPC6
tj8CU1dbDgd3nRh4Pmquz50owXYr6nqU5X4jboQrcVyxul+vAUR151m4mJVIHpCk6izSTSRJi8Nq
MVcCfgePEvxPgvXjrjG2hf+IC7IbRCvqMoiBUiybcQu6Hl3MsOHHNIcOL/GMNNCndYvyL2T3PMSO
qmuZMxzkusGsIUQGFpU2WwbTNa8JKzrrgmeMy/6gxvKqvnB3hzfUaDfDeGhTnvxH/5BUzK3HHmyu
WmXXve4lq/WU88tuXmy3xTTxtt3VAcHoZvAPkUUDUbwCgReB8RC+78rC6LVko2K8mQUl+OTVgg68
VM5lONwp5iajSR0G8RqFnruPRAKsabDGYkrLx5dNV9H72aZSMERShoZcIQ+8O8ssB9rEoA3Dr9Dt
OegJB+z/IkiHIWv2hLHoLSNxtFy630BxUuMW54sT2juXGxnkwfhxjqL2gBAMTsZIraoJVx15F4wt
uNht/OtZJ5Gtqh9vp8dASG1rlrfO45ayqZNKIQ7YWSsdz49kcHxYEd6rIa7qaPRy4ek3ZisnR3hS
pwINl5kdlYJ5GWvzr8aZsCRqCPlW6CcqKu7OkkF9Ol/OF+xjl4f30WEznDe1ASkXh+oTfCLB7wGY
pKh6u0dIArUyljYr8DEH+/JVCUBSMlBkLzgcz0N0ujrYo5Pu099XLpcMPw5SZdHKK8WL+7oE4GjO
CBVwx77khMaafejJBdcSpr7+kVJ5cL9RFLBEvK7pLBJ1MPcxtHkKobDAShrYFjsmRtZ6Z/ubqJDQ
8+/19Ji5QLjdbRBjPL70jq6Gl+59kamsr/R0Z5t2ds9e7+/hOCPYXBb7D0NgOryLUzr/10iu7dwi
sr6ALvVaMtEZmN50fBXVYrIzZodVPqo6i2/iE9PTgVGE4/OJzWgW54BLlf+7V+Qn1dLNdVqzGz/e
d2GO7QP9Wi050cuUoeXNIC8MZ/87sjQFK7ABleDpnFQiJ0HZtMnMXq/X+PEom/Y1Eu1PldhTkCmB
e3QkVymWhKXfu1mw0OYj6oXWeJ3zr5oHC0BcmKsu7TRDo1ECLIJEtmZB5T21jci0PePBLYtcSyf4
CAxnOYQriJmI/eqN7fxLzVoz7h7bKlxXvkL1vNrianGoZDl1uNjjK2zZbRTLJupz1urMAlxeHXxm
zZUzqKlO23MPTezKO1/Cry54qfLrEAG80CMs3cfCMhBDTVG37RcyIWR4ICP3FO0/2UYR+50PBSRs
0MJeAL15UuhIezdjfl9+vB6uHQfGfMd2qjAnmlg/J64QKhaDrwVo2erRRIBgaQuWl5Ki6nx/r7Ms
iKNqdosBcRbZd7Xed8gxIZc7hKEoy3enQMYD0o9aVK3Z5L1PUVuTlmJ8v3j6g9HbXkfjgQtF4dFk
EuPxByBWNlHWkGNada3pmV5TbpVvWY0uV2RjTTDc7cBHI3ZbXKMrSJBEaIhMZZMrBh8oSz93CUWa
HVOs0h00YP7fgKymFfVW/hKbwkW+bDcv8iG5y6b4dE1LNoZIhBvcvjUVG5xheKpyqk9CrsR16HZ8
8FdheG7bpkGx0UZ/6OTcWa6znQRhq+y3W4XV20KhFHzCYSFL94dFU5PNHlHdZ48fMsZBTBAOe9aw
RsG+nOpiP5vfmCqU8fFgemT/R6okCsSVmN9joaqus2SB9IwWc3zOp/FTjqdkQmaVyzCIRk+mrsYD
vkbH/2QQsmC13e3cLn7PGb3Y41XoVVCTXVTsI96nhjYJLPvckWQavP2m11GhmUL82VePS/7rmd4l
DQlFCftChZywIrV6N5pyKJ5aRPPAMCvHYZVsMkeBUJJv8WbZcEXobBlYN3KccjNVY1uBK40JnsBA
L2Bz07HTHGtY5WeagK5kYpkJqgbSsv9+p7wGc0YyKUIOOWHWC9T7nevQynHquq6IMfSpt1E2eIQR
BNmntj4mTJbukTThI5Zl5q8J5H8l4uVUgcDg8RcHzwwVapc86AjF6YGSh+H8MsXVFzHMx3Bixm11
JMzC4tv3aT6E1axTkyYrSAz84OpIFnkHP9uPeUYziChJNOTa/bDQcVzw0S6IKznLOn1B8BclpCtN
YU/lLGaOHaomqZEwpcwJiaZV3cLxnUIXStXPGkRBvgb9MowixuP3aR4KYt+/kei1YGXLxTCbfsNz
aoPoW+bisoA3JUXzrplpf7C0vU25UEincd2z4vRNn27xwRv3qjw5bVdofhWJ8rwbfJUmoXpZj6Wq
feE+K6lbG43kWMzO6rEdqpP6hxL7Tn1lsTanRodwiq9NCttk1yAjLEB3pTGWcCfOxOfALu9+ee8Y
uES+Q761wUv6JT8sE1d4azuLescstXKikugQPdN6wrYfcBE/Z3BvmC/DUgCXxWqyrM+3PKRPkgfy
eH6B/IkkqaJR56FOMXN4rwjAfd+UkvMd22XmsJbA/kqNvVFU0jypBNnYAdu+R7tXDKWhycRhS668
OrzO37erAz1QlYev8wyqljs7cyTXZSBr+YpSoDfGl4ouO+FgedU2lfwQoJJ+AZGn5JMb/EoG4syP
ZCv852KL3B6Ahkgne2ZqMjRFIvU26FnjLLuUa3jANUA+VDcZhphK/51O6hr0ZIvZLtkMCO9iNzIZ
VEjfPdI4trKJHDLKiYoMOdCuLHHRJEFm18pjvS4kyt2pgLPaB7jVLKdUeARb698RSDm5n7hiKs7s
jfkhOLKlpTREaln+siDzeATmC+7x1a+QeXfmTjDP+xmbrIuuwUZrr9O/8Q/kv3+JUwCZ+EQ+uc1z
7dnI+Yv8j2fVnrNC69hrBeK9AWTaRSCutZg8/K4HF9pmWR+HgRKYwAjisccaCTfpBtuI1CAx7S6X
BUbx5XddoAPcontURpInOZjO75yLBAMogIpQcMerc/5/nCfZ25Ze7ujnZBdxOTJtdaOKBuNL2Eww
OJ/VtJ5Bvq3AoTNR3iUZnXntf+37fUnN2qzvOucIVT0ouDWBaQYCtanf1flO1hz2l3uk8LxT/ubE
awwgVUkrnhOvCdTXI0qxADk7Y4SbKiwE2qlS0LmztussnyHmEk6SISQr0fkcXylahaHn2/xOnwK7
I2CEagyQ865pukSchnhFdfqj9cwklrW2I/PWif5gct15eyGAtFEfLLJ91OOz/b3tRClDlKu2F2Fo
iqXwRhCSkijQYdGl1IF4VRI0a82dkpKkkoW5xBWv1DVb0UnTIDK5X4J5Z2yj8HNBLLc8ETNziTSY
lqwUsF2OIuBQDwP4m0eKDXnRynF+UdlvqU0KfmyaNuJHsomipBKW6+q2Al30SNchfaEYLtexzths
YWV8V5XjygeYzxAM/XJk11wWYlFCOXSYPhjg9JlhFAglXSjchbzZEPU0nNNn0+IzVRpGviAUOKWl
9J6OoISKmuYlfyTvX07sGFvlbZke1W3MiHbrSAKHlq8CBHbbinuKC9NDEQV7FtUW2SUz3Nk0pjFR
AlDUy0PaMm4XCWC1NAwlSlrd+XsrSdD55PcyEFKCeUOdDdbUfKprtaE7Nlf6NF0OBUS26UXI9nqL
PLtUVJ0HNGi6JPZSlnxDjVe/0vaujQQN2nd8xIWDK1ap+Uz0Q3UdRKIiKEptUnzaSOfDY34y4kxl
8YtbIR1MImSGZARL8yDklfRmoK5+Po3pRDINBDX1xl5nFzlD57hIJZKbwiyoMlbsMbavPNgwCFFu
2vXORcrI6xIICMawb/l41UN9mpt4fX1Ftk9t5JuRdHjtqFV3B8bWB0sZNb2up4A2fLgwOWtNsuKO
klYPgwBLs5iDwg0sjyK5nT71bILJNJFycM1+Vfntpi7ADfXa5fX09RgKGBh3VH8sjwKWzPXfqVpU
0i05n0zXOM/tWZ39mHGyWOF/9f6ebvHIyKesxQU33TUcH1U/JY4tFuZCVdtg3D/pMw49I4MCWEQz
/4knalEY5mjNXxPs6WNuGhUAZ6/CvtseoTpV5i6d+eKBxB5ncVffoSKhTPYtwezp0I5+fSXksxoP
xVQ4riI7X1bsQWhwuGD1jYlTUnSBl1nY0VSyD9oq1pCClBOu4X8KdrfAllT0hAvY54RU1V469YS3
J4BK/Arbxzz0rpp0V0KQwA0Ve8DxerfOd+YbOK/x4OlB2gQI4oUwudZI9SKR1OG8gxlx8k8QFmZE
uDnAzxTBE6b76Al79ppTngboXAtAvi56vz7iXl8eOZhbArHDo8+AYPiKMGbl19/Zyb5eZQTweU95
bmsMtKPa9XmHFghTpFjvmlVaIcxDs5asAwPkbTvDjE3lBpxHD+BGi6fwCNXDzPo+YU/X2IL91uNG
+tO44ewxWJw3Robw4owCwHBw/RtSXH1MgmHeYfUS/xRt8u39aW7s/7JUecDu+gYBTD3ldDctnPTe
cWuN+AoE94h7SiQEDrEyBtGnUCxMwFmJEtB+VbGBhZT6yB9lIi+VlqDkCA0rddft5AzvMZ3S1qoJ
TJvDbk4lgs2CsnlHj/G93YjXlaqH7R6EdyJp6BXKYSDLCe4wAxPWHSI1TE0+oE5+oizFs8WE3gAI
rQFrtX7inGxWl0J+RRvm8S4g2Be0HNQ4rp7eOBQJsbQELDBhbL8/Kh6uTEWEOD7RQj+9pn64mCB+
V/tCWfrZE25+U7IR2rx9rGKzpXkW6e6CG8IuG3XO/xuI147kWzY5SoLnTXLfYWlQJMd0J0WTGFUB
vlUgZmmHghKd7Jjmx0SbW8aeCxiGuZ1mJtusWWmVOneTi+/WFomvqZ9/7VnTrYHDtQcjDBxfmyQG
N+AfJL14FuhR+3sFbW4Mk/bvyEnNLfxnT9HynyGDyyxBjnbUNVMc/S+Y1koiuYqPN1Eqs/izLik5
vnmEEIcTFtBKe/f+xAHpVcBTr6oCuIRgLrD1tVMlQ4uqkUtaDkyGKEMiBFlMaz7hD7JglLIXZnLf
NPQL6j3m2MyrwDZ7MWE4HtXn8GbVQnyYYIAWwYIqmUaVeHu/ENNabq2M8ktnEid8mg0GVmW55mfP
PfJ07Qt4v2+wvb6LZ/B/TZQbrj+q+/WkH+LKKEA8mzRAwJZHjvZGYhE/icJIBaIJ+I6cHHfbW6Lm
Fz7Tejmca9PhPiJ5JZABQjFHJ4MWB8iOGgtsCw5zJAit95fuR5qCCfrwMGL2Ka0jdzQIQMbyIBzv
GIyNvFskwZr5f3Ukg5UKgp6ij+Uyv0m3jI9IT7LI5d0VICSwP8zDuorgSlIX3TQWzkN/ctPsP90X
DYkctWBouGnvTBVp98a/rPmDGwEWmWkFV6H+SDGezeMS22uFQrSd1xf+DF3ufH09JPJq/hdVPoVZ
eow1ZYFArvki9YPR4s3m/tmCEJueD+I7lF8gYCRw7Z+5ddD15oM22saur4C1PH/CifBpzlKAKuIv
0o9ZrCRmokvFv4Ppc++BSUEAI+JX5k664RmSrQlaZ5qjslNm1K7GSF/bu7XJKZhEOqbsexyV5Bvf
nP6YkCtirqiO/7qh+E8gILS8YTnC7Ti6BR/9P3sVe80Qpu7beCF2P4srsVX+i3t01YLiB8qm8KaV
VBPCIdjymAXsWp3w9CfBtYTa4rqdcET+iwcqR+XHV0HnITSvjS5YI4dl8FmhAN3no4rloLy9o6dn
5QeT2/9lkgH9iJNLuPMRsqDRep/69mKW3VdjFTiHSClKfkam4ZhNeJcUnXOYsI6GxXcEVgs0d7Yi
XYVLeAe5ZQusJXtUhyAMfm27DY0B8FcVi6XUQJPZZdM9IeHikFxbaxgOR/2ybXntdEtpHabiweQ2
Il26yIorTQzt6SkOaOt6Zy068M5UNSY1s7p4P7I/SljujCuOeWn+qoCNSDoqsC/nS5F/h7ZLVB0x
KiOc9HyUEB0ro+kzIkEaxoCS2dvoMV1KfGnFXJ7h/8a02+Hfrf5f6vOsw7/R9q4ifo0inNfyjyAx
NdUcGEJOOVB2CIVr0d5Qm7XpvcA37N+3GQHYbVFjFZiWwGHCX2ojxwmg9LSJOGamvfSwXv6+w3VB
eRhodiYcoR3RhBkvPQblrnS3+5HdSmoDC4cHh75FP17uLV2j3onls+SglAszGzAGvjxFwoiXqimP
HY4enp+gGLfbRPmkTiCl2diUzsu+NIODB2LfIReAIi+et9i0PhmLZdHhsfzrRtEGHDZZFU2b4EVR
3VlvoWRATV8/Q5DTyfR+HR65+c0ekxokovWy9zRK7+/YwY/a8x7V3la7qKJX1gv63g2k2zjnUWMB
Er7gIKyVRJakLB6Gd/XXJxzez3BNmoc/jqQlR1D+TQcZoEP8rUGsZwrNBWMReY2qRa8wzPNA1S+4
+2O9HtAxbLwYoqXLxecBqDvrr4ve17sRsaOTmVmwRUYTvliBpY2X+A1oZ+Ji7uI7yB34gKj+Zflc
woGw6dnPkvOgQ6CB8H+TT+0b5N2UdM9hFVFMBg6TszxIx68SLdyOtEIlZ4QqKeTjIEnxuVcDCtzF
7efs+sGEoC7sV3IYFgoSVmmhn+0gOxTv/OsuvIIiqVQCcupud7nhywIp5xjBwHrDSNaHYP+6xMu8
LyHOXcyM9U8IpfIJEJT5GI4tctBX187Yr1Utx7RepDseXwfVy7ZOkNIOTGYNS6ahBG5DOLNrulhS
ydMx9qT66tBN3ymzXqI3jpZRkdEMWv0Uj0yzSUoPy32hcryi+RHsTU78jC9r+5UiT04RC1/Ie/kp
ql3E6phPecBR7JrG+ki6IRk0rLw/RiADsYHbRFCJ7maLcBBRZF0P+ny6phGvsFucJejYhi24y0JQ
x5QUbd70NiWiJEuCmtdL7BYMI22B45MB+ANSLu1geXjz4CBbq39hyZScJm71O9EudnaNNU+zefjf
ghFLsbMSSI+kWt2JG2slf60t97yyQjRZyhLX20bP4K1N12gNUsnSSBhkgLWeLZB4uXhVcVF2TUC4
mULKTqQ3fz8di9gNs/P/QL2gI2igCU51hHUs4Fx5+Qa6lu+GQkDoyOvhWeQk8WWl30leTqUi2Z1J
exHZWRBm83IQPnsd4WY1/A9PHj2xNjx0ID7Sctt6vl8pgb8SXazNDrI3UAvuIuClfULWqbec+y+Z
vEd6Z5ai2M0aFIgBRGiEkXSzUcWziCplk3KAdgiz//IuGALfQ8vQ5dzkX2gNAMl0rTcqJHq/xWl/
N9hqzcf2jO3s0J1lGDENfWWy7C0ppiqUpU9YLEAzsBvnqyEKOu2q9GbbG98hth/zSDjn22km7y8O
s4Csbg4XBvKEps6Ke7eDUSvZ0jWGNdN2CDLUKOQS92cZGBWVZqWwbE8FjrOLNAdPVFVZkGKrV7BM
ONplBMuHxCDv1nl5AoPRUzsY1j84fqCA395/koeLzKVQyGKudc18/AosgpDSD6PvV+FyK87Guqfc
wnCf9OBhmDayocqLlj4KmkjW4vszW6UrCQZ/Lu7arU9h41eUwKC6kQGki56jduJjjQB+Nt+3kmtg
KJaWDVQs1A21cUiYJq/x5X/DEa0aliVjiwKAjUwDPHYi+vIO94eOa4Vw/a4DnPw/IDyM1b5HBk9G
GCqjUnjjYR5QwypbFvyW7A0pX8L7PS9nhcvDpsk9WFZVsSccITEiTdIyYYbFOVX7FO1GGUl2eisJ
JTXuwHsYusQwhOZc/DAK1To8/eH5KlEHRzGgJS1v/+2nfxLGDsQWLF/iseptGx1xSuno6HD/8b/P
D9u5hHaELFQloFUx143ce2BEqKnArKRF2nGSu5minaK5qNw8bfnR/PNoLr6FbuRT/MnQPVYqKfef
QfwqVLbUg8ULosuresAjtnPc3Ug+/2WgJkvNQd0tVOlmxqgmTPp634cyaWABm3uLMPG6fHrJH8+6
rsqNfB2Npt05AoSfkTJqAlzHoJTXUDnIgxf/1QAkbHWbzuCAEdRSmgWtK8+gdG+g0dX2slIr1Ym5
9Y26bidXy9/4TwLqatd7C7VVYRkdhJ4GmxGBHxUWFE4hyvey/RqAWjoh/YBqiIlACBGJNKAOEYBp
vXT9tuju6TDBJBehtr4Vu7CcPpSFKFRnnkvDfxj9ftJrQxG5gPtqUfVCur5IH1J79y0h1GHoetzF
nqM5wRKS5AxJ8AIiBsl09v5ddJZBpTpJymql2TbN8p2XR+gMmczC3qn0XjAc0ygX7IGjuP0GARyQ
xaOGVGY6WMwR+xs7A5CUWB5KksEsQ9eHBmhQE2JimM69XjDNz48VUkEKZZa59LnV5mSX9mVZakdq
TVdiOQXBUbjAE3WE+AJYxgk0wGyyWu7RYTMlIuPyJuu1+3osPQbp9NgD2kvXvxRu9kb7kb8zqO7r
9f3Td1n6MuTYaeR6bgjbbYfWA+aBcFiH0ruLL1Kl5kfepAOAPRiWyHai6KcNkrkxbJwZ5MwiGBqr
aPazsPA1Zrka/QDhQNn87R3CSccyyF5SE8p1WM4Wc9WBHf9pS0HHPTGg6aoJsij9Qntwl7HtgkrK
scTmEOo7J20rGUDNNzmBd7t15tk1z3Dzc/keU1/qSZ7AhCON6xP+yypZiFJa2O1aDorzbTvWgasw
lfIm+SwhILN4GMhJ/k/Yg/BnDW36KliJdd8NA3+5ikadUDz4V3BhKidhZIAfXVMJpvCy2eNA4IXq
eFXtF3adWC5RHwIy+UM2jhd5DbUPLHfswhkvDWJaGoI/JNpH7lJZz3IVOJCrfOR8ZCXwvUXowh2k
LKIN5TCA9LkgP64mbgtV3X9YAXGuOtSNu+kgCvy9Qii76Bwz9SO+clRZmBOLOlR+XbptFqCwsDei
SYHviFh8gM6ZbEsZfg2CnbCMq7utVdwo2OSM01ExOdU8ZxNd4Cpevs48vhn97450R1BpRs0Q8BIB
XjtQRpeM0RO0Nw8ZK7xGsko3OeuMiK3MhgXwUJ2iqp+7U8Axq5d/lIDEC7+n38u+bMR1ZSccu5/U
3MxtLQGucg+kfmdDWPZ2fEeukMeeqmnLurzfFp9K4+0b6nH89Xhm39hQ6ZFQhVz6+wlWesjoEDKB
f2Yrmpb0doutNdmJk7pxSckoLbw0+mXDQ4o/6sxboq2q6JDHnJFYYqMTKvjLnelkdXe/RWW4APaV
jUu5yWqFr8DCJ3WvcZYfTf/mg2rbr3h/+CUnZWsyWVxRNcmdwWE3qcxQ4yepo61wmdqo28U4m1Nv
XUQlUALDWtbWYD8/5HRZPzq1cgzw9oacj1/PlhEusGXHUieVKrQHFh5OW7quuYRUErZ2Fn0u3Cj0
CWJMCrNgqTMjUzht8F2sWEBRdGjFQeHGYw/ptXs0EKEZk7OZwLXNntfj5UT7O4L8/ZE0z6qM35eB
rTG5BIbgNkJHi1nSxhghIZhTlOoAL0FFEdjGsPXFWhj5mioq996UljEH+GY5qu1T+NyAgnV9C/kB
ucIYr8chTZV4+xnFs6kl9tNKkUAEiFMzL8SJ/8oPt4r/k2nBEAaQdyukBn5y8LQHihKGDE7LO8ZT
g0wZuA83koHhr7WVUWLwUFrLGxr1Ex+cAlF3vcmcjVeQr/3yvuyycL/8t2TBUOQpVssSQh6jsIms
yww92JRp99AUlv3Ne54A4i0iBHyTvsALNeKI6+NRWxww/YEzHoAQk4ZSR7BVgpqBo+H9cIpn5Kfp
mS3vzR9Z+W6Ks8g5KXA3jiOSMtnr017aiMaOx6pTp0Jr/qsACRh1n1DD4av5YVEbHWmfcNmd9ppl
HsQVmNZO6ZlifMWTNgSVueDXVUbKjmaNIUpGUoxvzu2Dzy/8Cau/Y8yi+Sa7nkYI66JWiePlM0S2
bA+eJiRY5/DLYmGKoTDwH6W9QN711bnKBDZbRCspLSbqIGhiUzx0pBCaxqLjtNqStNvOP/zZnBEk
Tiw/hMuyiGUrBziQ6v6dWc7SvZR3DQOMfQ3FkbnKYoiUzEp4l1qwKPO3GzDx9ODXNks8nO7Wy9sU
Mxnuh7sniVgxEFe1Cn/O8RT8Qteq4K/WZaZCtmnT1kvP+llSvirhIHaJMyhh6YgGrLR79yUfbLjl
5yq9jtPjfciTPpJyXrMJzBgzUi8CSSSjf69DSkTe6rn33OudjTbXSKgbKo/uQckQcJOISVNewVSp
woEMPDHF0KiaTEnpnkeJ4HvZBnhXc6gIojvXvd3yyIoZfyAHPF0fWQt5D/xazbK8CcmHSVNeO/DP
81bPuQQeT0tVQ2/MJfkAymreRuE/pxfc5a6XlbRvF80XYlD/hbPQMkFmBQjmslACf6A58/ZQ4RFr
mAoJ8NIwd+OYSn5Cc6eObhoh6/z612w471+qUuU06PKYnGaPti4Xh7rLLBK3M5vAvuYeKGU0YsHR
smmojgr9bCvifCs+L9vBW0cEnQumdamsa4A7MHg51Jd0J1pZ6MGwjCpFhWXlRTqozlFFTseChHWe
x0zQARfvehvd5ES0Nl17FWBC8lExSGCXWpdbE2ad14snVthwB5wmv47bN3uUvWNrtZpIpbg3S23G
jZJI41Xy4TJsl/xjR25jyAzbebVVf7/9TX9LjxZ0DreThIv1JSnwMgnJFyXXhS83a3fg0WxYVPaz
QOfg81Tevle6vS5qbva37iHJley4lM346VO/v41lP8defiBUT0p0Mq+Fjwxj00Jj6K29F1IQvIx9
mIDcDHu2+zNsMTkHCM0CuYkKoByEPKpziv65fOLHeS2claIckPXt0jyQxdkp90P3fLWjYsVUqjZg
5P4LMffHRNRVsc8BdXu0pQfvQTWZvNQ4+q5WlLibWJLsmlI/g0K3OkKiIUnqKzqUoghFfgCgVKaf
Xjuk2fmtTs9ifeqTq5We2TyScLQ/9TkcmbVJfNexq2cXQtXi0grSUSlpaDfZZ6ZeL3f6xya7ZAzp
D5JXwRaQAjP9leZGnwSLr30Zc3VuQGTbkVPLIECZXhDEniMZBmQrfo219HIktGQHz+8j1Q8kPUoM
+L7HdaHp1/dLM313/sniAUhwoOR8hdyGh35kVOIXadLJTRvkXqQDzBfe98iFhpUpH1nBEGka22tO
48Os2wNevMX1ihsRuuHeQ95o+WHhdg4YvRNfSCHiy9KzJKKW8n3tNryTyQlcWiOZCdcM9EihDEZj
gBSN8/TPmwti6BS5QiUMr8Rwj22Tas9ubeBNAKf/jYVor/cmj8Avc/r/KUuFQC94nZITV38N/2aC
h8ZZ/3E1j9rfmvVUHof2iWFY7j38iz0hiroSnwkDdlSXF7Bxq5EfLI/WiGkMYeupFOy82mYehN1V
LBr2myfZbFyV42B4WGww9CODeX6zXqYl7fvMh6CTCMYvHnePA1IKZMeg/pX4cgqW2JqlZk7mS7np
gbp5jf/ZovQVlh9tlAPnwYmoiAQw3ygycWlWA061HLSH9jAaeg69iSIkyXAl+FYJ1gZjTxRR8TOg
diz3fDkbUBfRk6wtcG+4K4Xm3l+3qX96utiwGBdMM5z0OIMc7w88uvkOr25tOln07hZjKxHYM9Zr
/bdDotHK5GP/sreNr7kCoYC+gRxfD58iM55MXN1/pk7R31cl0eAwDgw/zNTATHehS0ZujBUbdv+2
aeGXnZzX/tbPXc5R2NHrqEJJRFRIUAcSTE1MXTpcD10/MTjAm/yko7uqpg6zn4B7YHYpAXSf0xi/
T0cDkHMM25YwO42Ej8kJLPEL1MaSF2iLGjumT3XQZyQeZdo/yEqzmG9tmDbxPXj67PHyssoiEHBI
w4RbNuIxf21+3a3Yl2U+3zHnCr6RKGBcYhojhwGtKqxWovSJmQf3jHo7THpwdQv7551qJ63OzHgt
cODlO6MSFMzbpk42Ut9D/+UrrdmoVYJH8vOgx/6lUW+MbnvwCfvdFeoLyx7NEmxxuyEGxhx5o2c0
Ox6x66gX6hLPDJpdjYsuHDPEYMdm8rjwRtkuP7NBZc0Yp3vb2vgpxTrrXHId1T0giz0Gn3bBTwgp
uvtq6oi05yJoUqBaor/CDginnpqEHDNoEy+U2Kg5zeROOI9H9Oy+ZbLkyUqIOWQzc6QZIa+ts5/j
f6SW02SQOn5S5WnCJdyB8+Mtwouk5QYv0CoLfszFTM3G76rbvRU4Kuff2d6DSEyVNfOk1DfJU4NM
ERFSLqewPT7v44Hyi0UrwN6tg9mTI79EiHKKwUz1TyqDzLpJN5S7Uyc2u6wCyh+YRUmYrLVQ2Nvj
Ss7jWcM1JBDxmBaJb3LIv3qCT7TB54/Gtiny07NOEg4aSG/iIzfXZYqe+vkbrVM9oTErpF/dHMkw
9/Ci/1Cviu+kudYhlvHDDwPvNXEcp74EoEYMfs1MtOunSfNTFcoaPpbe31TaPtmPDiuhuYloGKln
zYRNfRbfztiPJq8BifbM5KOIFaBbjnfYEO/P5xNZLxEVd2nXuZgJbeLCscV5pm199DHWfpv6tuwt
hiha0IFIjxza51SxT6Ty1m+WCKj5wvUHyZHWGCIuFLBth1kPMC9+YkoUk/EO7KNxn1H+Vlxs5qua
5PUx7V65GxY89MhZxcwUvr5fkTbq28v6LqYO+80rnk78Gw+9EqXLJUFEw9iGL67U/cShr3SlO5i/
aTcfi9IR1TLupubFRW5KDNddwozoi/2ogakOXmw4QHBwr17am60YSM+HaO80ewEDhE2XshLQ1/ko
1wsZn5S3Bjdb84Y3xeJmCgXifG6ApSlMHiO0z5zAJRYhuOqDSVVk7xzC6MluKYL4QMIB6D63z8Dy
o9soYLdn9P3piwKVTSvT+1qWOy76pFhM1qrT9hqA/8kDpWqaEGH44hKIvFuhIOsJWpYFKmsqQJSA
TE8m7vYHNBTKYgSXg1q7K8GmyfO4IS/xVluEkKEGwF9kjGDiTu1Fz95FsW/0T5H4si2HsjdC8lTg
6TRnE99hPqkipbRQk5efPUK5WzpH8hY2ritk8gX1SQ10wQR8MpWsqg1aaG6s92P2qd/VRU1MXW1I
NLXsYSQx+d6zApPuIAxZnvPjkxsxSFoO5ezTcjG4spHe3be+4BhkSJ5RJlQwTZapuq7KFIv7SFTs
jm5Myi+wuwJHWvcxSsSCsf/hc6Km7KuKHrH9VNUr1dRsTyeRnyR8dJeooUkaTf7WDr4/Rgcw+lgd
8KWi7Jfu1BTFruHwQ0M9pHw2WH02UrCg5KOcLJH75x5BvYAtjQywjAwXvVCfd/MwEo2nFO7RlCoa
/YBRsGI/CP31dB82LtlgSPkLwuf8pmTgUMDyEtyqnS7pFKXj8ierejRg0hrk8qGRxD3KZ7QuTh9p
28YvGCte+f0LzhpqANBeCk8RFijKfoCuAwjmp+niRyWh+zDPB7qEgh7aUrMr5P2JA0EKwkhJYI/w
Qu2pAN2IfEvA2AxH1Tmb4wYjZcIuSlIujdIWDt283VQSUmbFAPN1CdbG4Pk0j0es9pxaytpTD0ES
1SeBmmam9zF+h03fRh0pY0QZXd2vtKLFTV/bzYtofU2n6KQmPBvuAQldNce+OaImUg9x8/hy1MBF
pFtmqJg6IPDzueK/0YiGjq15jClRYRho5h7I0BcpaQlRiubqtMLJDMazsuR8N04U6sXN7xGHWltF
DpuzNAR4T0oh19oyVBFGaYA3kP2i8cNCj+QGTBfvfK+rNNR1OwOJu0rZywZTfRuv1SE2pY8aHp5I
G2PoAC1FNtFapjnBRKo8H/3fNBdR8+zgeqOZ730L1UUsJS20n4A8Sv5Y65vAshJg1153BpipCEtA
h7Zrl1TZs/ASGkcq5UhNS1T3ah8nR5DKOt9YGxnEuNWLuFPLwoiSHiV98A3qxJOtYVIeXtZXeQiN
VYacvNbyVKTFa/vhaAhNBbEZReXr0lGACoaZnkzbWFo3tJsS2XMgeHoFSLd9Ku9CIt0oSx89M3q/
ZW6Z2tULepZfjFY+aO+TOSmVLQjiQYkMIgBxNrbARmlOVifd9nYEcMNhEmWZ12npGo5dIwI7Sxg1
G7FXlqNuBRijnDm1zp8eVjOlUod5XD1japSGTP+SVHvhjQe5qQhSdrZiXTBdE+tyD89xkQPlrV6Q
BOb/nLdnr3huIhj2SW/nV61PdOY/0XHwoWwcZ4Yu7mtgTr8a4NvRAd0o8VaAja9K6hbbfQ7dpkXc
9hLbx2j6+r+9ZgMpLFDljJAkZnY32WGUtUUcTH6+lHaOCtu6ENM5N8/7KzXuoiiWdeBwqchxowtV
Bk0rMfJIZb2shcXc+8DtLwrgFSarv6lyt/+/ZIiz3rRKu009NNhpZ7ffx5CWRCd86FO5ux3L4rNE
ekgQS2WoUAPhpCkqXNxeABKxMxjcz0BTsggKaxJsXMpWz/v2VPlKaPi/BzikkvSPndAb8eg+lIqo
vM4j6SxJ+cuTGdcHSGlRJ3cau2WzRKmFU1nbf3q17r1Q9e0xmUhlug7QGfgSMi5BHS60dN2OgTCR
wupDeji6UGKcr/d4akhg0Zbl81Rln5dV4gmWwwjH2jqEzLeUaZAimA2oHTsnXJYNgM/uWcIdtWzB
P8rBp8TuH7n140XwsdoZVjHqPdoAPqd2cD74IjDNHdTpT/Mj1tMwJA+zWSuO3h/CXXivYdLhd303
efCf2YbobVnn0laab8TleFalhw9/vyEl93aaa88nWECtJn11FnFATo6qbltgQd4mLjM66viDpogo
6wkKJH0D2CnKXXuv7tGB4g7rz5LoUSXHBIXuqaDBKXO4aOrAjvzOy1/SaqWUvHOonY+qjv9YsO+T
tW3cJRjy3IV2MbVBDl/8Xyxbk3GTVzmQy8cGK8r8Gy/Hg/qQBKwj01ssClhCgEB6RG4G+GnhM8Fe
Qbb1unjF6Qto+pBGIake7bf0uQAPqljgu3jIZFk+JjUyuUY/13QPm3N8NatHehxfH8TTiY4eZdZb
n5HoiWKAFonRq4uGvAwP8ifq6AKp5OU62WWniXUxdpBXMHXvpmtrQiWw1HQ125yk+7AXa+1KmCwf
ITRk3QBrmQB4dj+HAtHcQ7qo4d7YORzH7x+JfjdmsiwiRjbLKzamGGmU4gkjCCyW+C2ukqwVaDcZ
lvbUNABeMbMMMByf1Ss73lXX/YTFyx8uUTpot7A6cJiIBZEbJEtq8q9DB9Lq7ZguWMQqdp2ITDd+
g7SeButff1T/Jnu6hhQ5faCGuRK+Hqe4ipMBpsrqNkoR1hkG8ijot2B2CGr+g/trTG3OPwIiAZzI
vu89v9WHyUKs0z8VB8MshmBc1wbYZ3Qo/rKXWtz2lUcQUD/hmUO3RxnvhGjRMlSNaH48TuYztExy
1KGJNGQQ6nXnNaT7hxoMB4nGMdhELFipsqShN40sW0B8ykq9MKgRx053wic8RbeTnqS4ElzrUwxj
mmFbxCm3pzs2/tZCYc84+k+YBwv+wjyJZCJuXp1ZPbyKJeZvIzkXswpEud4efYcWRNDwkQBLZ4rE
XhLn5J9xJus4lvVvOSDSBRYfgOWHz/WWHH9dRtYZ2uCD4E68OhHjSSDhX78192BXZMOQF68ripYY
TZ+9kaoOV/UMzu/esVUFZjlmfOLB51Ka+Kq2o/R7YfN0+Sd9BY0xEMxU7wkCCEgor8AnLVZgZkWE
e6eWxiF3ytWh3uB86GZVbU9zvj3wInqvVJB/OYU5QvuL02pqG2uYogs6bTKtuhZzz1+pd3lEkZxt
1S5HEBbAXx1ye0YqrSMq1243Xn3SIHPmJK5y6gFeCND17zylXM465wcbAd7V9c/jEk03EpNuL6K0
GsfZM4M/HGoSoo1mi7n33tFjMxdNEc8Rl5iyiO4wFpbUMPRw3t03BAhpz/IvJdKgOZVB3bO8ReoT
aKweVoReXNub2vRif40HLUiZwmqWxr+ot78dWEr+NIZZLNiESEkgSR/PbNzYM9/SXAxWh2krbURa
YdKAUvwJ4F7XqXOhdU+zCEx5x5Ic9QLsunmaiW/6TcoKiJVzA+KphGCqorTPTJSjJEWz1ypU31eQ
kOy5jXUcJt4yx80hEdnjtnH8E9OtjfLpX1NnLcEInHIPN7lmYjR09vtfFglkvWR2PL4ld1AsK0Rj
oX3lIOyqvYQtb9cqkMb+X4Dq5/oEmow7gwtkN6RjwjNWs8JxqBxfwAzno4m109NxKVTZ41eUPW7M
eFKOu0RZwZogvr/YN/Ns2R9VdG+J2cvbOTNo/cwWYDn8i4T7iOVTBN7ZbT2ertMbrD3GTHbQajX0
DRy7zxE7bTdJVKAyDX9ISeRzPsCGlsVXPbEmDqsWM9Tf7aXfsU10rHXkoduAJv2lnLWXtEME4bvy
wV1oRqwn5cqKFwsoWFFKxYWBrzFEX0BKPYzKorBONSAdCu8HcMjLaFYIcXl91Rrc4ua0PmbBvAto
cVXZp9acfe2PZPhvm0kec4bSo0H1goMUFll91WJPxf7nlp6LQ38vAENw+hIny5FGraR48/HavlGf
kPePnNDED5+aJ7wzDKwjtCypIAl6NIBenqCPlucC1wRtiDnajuX/eMOU9ArbQC6pzyGiowjyE7VY
B1jjXzZQy7wCP29UP+DgsEm5C+CdTziytyueTL6rBu/aNlkNm9QlFv8MVEWVAZ05ohgBicci/DpK
IcLHRNbhWVUz9yAKgNweoTI/R4eL/4DdTtGwJn+gNsUg7wz1HuJyCNwO1RpNUdx03x41QIAeYF0k
1lilV6/LykoU68gLFiZMMbW6pBRrB2D6u4vqgdnfuN2967xeq7X+mct7V4f+l5OAYbqbJ8sq1CKg
BLjGOaVs6oyTk+mAnabNPmAgvBnykXfa3pB5BHGYAMHo4nNqQCyzlQOxijh9kHh8J1huahMqZ3Po
qYYxAVpjU5jfAWz+PtkcMUsfeWM3nmtMxNULVEupIOlKmlA/2KMueQw7m8maySb4fhb+LT2XfZ/Q
7y9F/Kpx54esrrpFydIU/sSjFG5PnbR3gMwr7tFYdVEV1Qk62QZz9paM1+Tj2S1k4KBM2RHDlzSe
rC6SIDyX4Xe4ZTeJYwosuBdwjExpeVELM6JiCGOANe6Ge7Dtn6z+Q9rpzPH/f/IamH9Khl5vgWIt
DW41x7rHk8xC4TXPX/1zpdNBzw+4GRgGIGyvQOxSDkBn2IYrb+9c0THWcB9g7retbsYi3rltUUVe
BG/Mmn64HS7L3ZXXascdf1sHxEs0Sn5CjHbzN32UB8KTdSOCAyM5MBhqYvtMOzxpBwyJ3Q4dQ1RJ
xE8TH/+w510J3bjp6Z1Uy+0lx5+WbkKscuUhA+2EY/jv9Rt0Me1KHEJsTBqt2wp2GLowGSR4DHKM
NhMCkScm/HnbMnaG+EJRkNVX2yp4sPXazacBG3uxd4Qz1Dp9qHCcFFGBLJpzUDop0fWZDDhZtEnj
5GbuzNjFgI4Pe/BZe/h98G2sY8Di2ERmgZH7IoQK+YxmlLX43rCvH+ryyFxAJQZ61iyAufx/16+O
hRvjmXp0qOoLOIgWjcAlAEjCPSB54FRBjumuqFdvgmTUMNDxxLtX6m52rsH5EAWW+O6LcAECg1BN
bhzmugJBit+yv+43XFI7Swqb4pv6GMVc6i9OqLcGYbd0MzOpdU5MNp5LcRfZrLWTzmk4ZFJ2pSo/
eaOM6Yv3OGk5HJMhJD/Yb+3kIFwz62/vrQ6PfiRZndnYzDrveWjfJWHp2OrhSdRJXdNlGGvWRIdt
z2UgbtV0F1GBKwIqt6uBAPZvIHuv/4PPBOzhvJi6svRl9+T4qdpXfSTf9avzqqgJHxbSRPLjHFHu
ugrmgAh2bKa58QB7d0bHLzBDDdY8oF0eHIFtVIj2qnlSy3bHpi6hYXKAstRCMG+afwIQ9dc4/y2K
fWEMO/lOTY0mzVfVRmnbBQRjPyz+hk2IKz1HSLH7fSkptxRgve/rksLAW+jFoDwKFwc/pw86jR/E
jVtP7rRsY23lVxrUg0m3FuOlA/xiZWmhedkL6ts6mWF7RWSwR26ZbJy1EAmnhsrIIWz9cOrV03Ql
BVijhgs4gam3PHLecZoqBNXgoavm1Oin19JSBNV2Hw8H9fbVWm061/45xt/n4akyelE0QhNBbM5m
Ld2qSfLh0DcUdkN+3uA5JEFcqkVTmqUa0tGdB5IzYd+k69jT+JNHnXZIiYz7WS1DI0RsIjJXlX4W
+xEDAJ7cPQAvask5myCT2fgSsUeyFEn3UZgS4mDUyISgila2dGy5p8SD+14X8vWxmgnPLwzhkKPE
Sck1Vu7JX2xsq5fCSagrgdWtpkllgZ2fHRTVyGg2amI6YRSYdH6rYosDH6DX6hXeuX5xFOij3XA4
oEvdcNCrWki6TaZr9zEzOXnhoeAynthm/Mg5FCTwn7w5dW2wsXEBjNwFpeCYqqtqcfTihHpO8qhA
Hc+hS4sP/fxMOOIYXe4tzKZPXH+c0br6QDmcry0GuHAu8RYEoAv/jsA5UVuaVMdS/58nv9Hra6gj
9Sw+4D1rBZOe7uaouRBe7otcivclBNm+egU3GubHPX9tl4QT/QHflwCOG5keQT2z2/yXoqUT5wIk
3udiwaNDfZlppNtQLUrYj9wsc10fMRTBlgFlK6x7Nn9L0ZoKU5eglfXKtaNKKX8Qr1HyLSzCqk/X
30hs4j2xCuqxO45t9kwdH2scFmIzNBrwaySOuDsuWnXr4viRiI7dyWRKlKySxa8guj38nuzae1wu
succhW+0Z7J89fOJ/yyKfy344rc8Dvs4YZOxdUBcocipl+cWcHhOL3nf9wBiyQT7qOdpvyDsr56E
aXcrF/xWsPckOV4Gew9EO/rR8RbbiFkwp8lg0cGMj+ItF6Ni+l6QNXynlFecWv1iTi3ZLZRkf/fr
dMR3dAq4czsqGNptDz4ve6USp2ZIXQH3AOCTWxOD8PxbY5sBBv+xTMCeM6wH8OV4QVFCicuR594s
RtvoD4nK+pdOKMdtj9j2XHWGXghyMCjjVvQmcciMWYthNQ1La7oGxNsbIM0Lh3Shzg7kiCWnVKh4
DixhFRb+9OOIany1L4xRfLxrvemRa5j8c73oEsF8uoFUZ+QBHNcopIc4VcC/z40KAY4+KVRfA0UP
ZlUFnF2sMqIfSK/zzXgDeIUa23UxRV7ytT+v67DYZad/FF/R6tpf5xR1iWIh1MZ/maMzIFcf9HYP
JdlGU6oV35bKKwetAo3vvjyPXIeNIOyXCtc6CisE+MCbgS4fLtErKXGNl39yPypzL+g+O71F8M4z
JoXrNEZWIvsvimKi3RV+OJ6CSde2oDJJr/yzl6a8YhChh1N1in/FpNSuHn1ru+krNgAC/P+q5awM
7O3xtOyNXdt8hpn3CvHCAMUkkuqTc7kZPQtSsSR26RFK0ruUuvofxpHfWjYhrU455RcnFOteKLcZ
fY+y32EntZhzNcAsHBUH851jWh4HU/N45R5dWBzKIW5LV6sYDPvK6DL3qVORfxa3T7cu0jCO8O7S
BL7hAD5EeYAAcTNAXtCWFZx4iCwMrJQVcHJznJeHrTMzFVF9G9Qw5F7OC3JI4FLYa1Qedk6YdkFJ
/uO6dzbwEm3PJDvvVj12x1c5XNHB6ET3qjoXUic627zt7Dm3t3SMvCX8ksEaJa3+bOYPpBub3l0o
VM58AdT7KoPiEErBOC8QppZth4NiFCUWmpq+3kzgJFVp6vbaxvQgM7oG7wGj+sPefQx+WNYIdf3V
n1dX+HY8SSa/E7o7TQK7aQLp8OxeQAKImIV80B9Dye0mAdToc2gHcOUDVuD4FGaMTXR0gN/0oEQw
1qZPHnXrRXklIAUI/ar+ueSsnvMjeDg7klQvUWuSFwWfFlaIGFf5TKHtmG+IpmcgtoMbKRHJo4bG
6aOwCC83HUxb4NBvZ8PTsacDuODWXpDZwb+5cIwCEwuJYTmdl4pF1YkScbZQHSs7FPwknFc+ln25
XzIiW6vkt7oJHByw74d1HCrgw53xzldmHCi81FWNdVatUi392Zj7hYlstpVrSNlEd6TS1Iv2IfD5
x7H/XZ3VoqigtguRNnE3qYqlXNWspz7s9Ee7+VxyGlIxwgMGXvOKWDegYbHdC6Z9RgszNyRJy3q/
5EMhKFrb4JQAw5UFx6tiD0p0HA885JHibWwx6zBM/D4ZeF95jXa2d5QbchcBfXTMNWNrG6kG97vZ
1vj3il2aBs202n0SjK05c2cqOHXnnQhutSNsoDAsX7Wz9BPdxks0nZuf0RTxw2nMCpov6xVEt0xh
5TqpObEOr0dYfDKfD0qE9jbnZQsIMkSBL4I52C+fADFXFPUctUTXz2WMl3dE2Mw9PpCymSxV5gBf
dR1fdqXkvuZH63yB17lbBNEhwzW2oi13GURQj/wbfOzCLF1MdpHdAmzKikZ5R+Y3/C4EfpxrGEMd
21R2e81gfyAQEMfJzr1VFgL9n1E6hQY5qYdQxMzYHAzK93C8OaTeaysAc8YvDTOMtW1SgjSW6U6F
SDPFjBWgAGVrQByWjyDOsyXyeu16Db/h6yjOyuXHOjAuEcfbtp/V7bgmIEYL0uOTHrN3IGZuIvdd
U2OEG9wx+FWv+4vDm23bbE3pqdjDPwWj7KTUB+7IGfcQXJ5/jHx+peELeR6C9eINLZgLV3shhArs
oFihoGGxK/Y69NR024XwYClGlwXQHysIeZu6nqxnIxm9llQvQLAiIl2O7H8hz9KUWc4tSRm1U55V
N8cmspNKcL7RnY1Iurw0+5Degt9QqXa8nlOymoFA9BSmGGCzIwYj3g/qCq3F+UfHDilruLn17Jk3
TY77sX5FT0JVNhcI+jJiaGItBvsnMU4bl2j5fUXUZO5i58e0YQJ8S9evvSjWuB00VvdZ2nhRIohN
eh6SC/kEdhuFMpbyolKKP0kAmC+s2oG5X3Rlk9Hti1fxcnCh+1+9XnO+NqtFNdaR0OZVdhHBynAc
sqd7pX6mkCFkxZ0argQxuAFweRIsBtThC2szmCq3a4Ij0PLvrENtJZpi4msgtW8+ccmKn7BgVn+u
P+4QCMlOqV5SKOQSljDHLcOb65r1MdL5f9l0no9O7g2TppFq4O/sV2KIB2cflSmPPV2+nISvelGm
ue60Uniue7hwnAhvSyXAM02iVzNhn3DkUo01JXdPCimyy4wdJtT9laBtrpwBPElF8A2Jj4zQ/vJw
Ta3557o9zPJ76r8Fi48vF46efswVkMqq2TZGrW04CJTOxaE6iQr/vCVvRWrAfl25/nn+vQuXYHHP
zcAB5z5QtxbUj73BRUtamfsrhnwSCVd1poLMZcCYFHHen/QCix0qJHL0ZY8f05wKUfpkeVjqr6YP
zB61RewS2BfRWTK3sOFY9jqbLcWkDnBZFkKZTEn88Oh4XAxz/TXue8OzU4xQafHLxIrRJOEaY31F
l+X9VNB6HGLf7QLNNYhiotiow+UsDHqjAwYTID6YiHYDFZoeIUfmTjvEKB2W7QfVFeEBB5BT+xAv
WaQ5yzmVQdr/XPqEuKU0B3MOi8+lra2jOik7kcrzYtZPxvRATWuuX/myCh87wjnFl4LBzYlFWYS+
kzSKZ8H/JAiiEyKtwybmeOHjYoFK593B4SFliEP45YMvmgXwmM542JbbIIeOjp/l3GXGBt3wUcW9
HqmfwODMIVf9ZeqVs1Xe8O+mbJ4AClqkCnI9Dmm0sjWkYRjxBre3e3yx1ioWKrrQE1/vTfBuHM49
mOux+L/LXkcyRDl6+DFRvtDPZXC+v3RlpsxoXvH3RUqIYHoFjWyCNALoopsc0ggYi4++vLFMGV/x
DgvbA4X2y+eu1OxgvbQzMKrnnQ6FtAblzmE2/MAPTzyYIJjPVDuQpOC7d96tY5m2vJJJf7KGfpF1
QunBcRo+LJCdHpjeEFGPbFsJaosLCCC41xO8YC/jr2zt+fv0Tw+/2mMvBlIU6eGgK/EpSnFlLoHr
j2wLpgg3zEC1p7OP2u2vaEL9Sak1EFfpGhloCnzGMYdCVoDCesK18Kt8Ii4u4rHpp9Q5exGIacYq
baHrnU7OxTiAIt4m4BFNo/9l7PZE1hZRnP5dtoTD3lG25OBuMTB+mwCwHdKoiXS8V7ikuPGMq5BY
vBLDMxWws91lLl96I9i5XTUX3Uf2hU6ds8fIbb2Sz3cUCRzFNumXH6FlUGpzpMZ6uNIWO3IT5QEB
+qqc4I1Qc+SJ4tU2GfVbtQLmgSBUNDnaOP1btLlZWkGnDTaI12tM9iEY5I63+NH18rJsiK/iSPgF
NB2H+SYVAw/DTf4/tOnaemV+2XbUmiPiGYXUKFBnWNHgya3efaYeN15NJVkr5Y8jEG9JPgjqU4Mc
+DI82AlKTwLP/Gfv/IGqMBr3+Kp+SvumvXHnlMUHzgFTE2y8oQJe/9CUtTK4OPTs7Eyn2GW7niFo
zufIanwYYAoTVupJ8U7qB8MVAiO6FMbIe3Tx7R1diVFms8TG6OguIlfkXAJ8TLHNjTil+SUxSk6X
9XT6vIT+luz0I46MaeHjqePoLHo52NUIcMAfebn/+3w1KbAmRN5K/3m5kcNG52ylLQV0FxJy/Jz+
Be5jZVN51wLfQmdSzIwd1D7VDRSAGAdnRtDPs8ABb3JxM9Kn4NPMI/mCnMS8Lv11iAkZfW/u2rKz
t3R+mz2tEshaepiGdpsx65B1VDDg2GsUO+BZNZXAUU5N90gKCpMgmq56UJCpbVzXT4uy2oq9XXmf
jA0JTHzDYyCnAr47SPmKN87o7ES5Iog+83TpOzxUUsCT5LOS3T1VMskv/8STE4E2SLYRzsfL0LUW
jDs5e0805p75B35GzEpN2HHTqp7HCC56WtgoLfA3pAHZOvO2gMVYp53LuoeTrFbTeyVwKi5OMq/m
Hijk5E8wdn+qEsyqR9e/1vlFuhzh2zgvfgqmFRLe8QZxVlZJ9e22Y+sUFS7jGpy2kWo+93juE8kb
epFUOOzE+knOlgPGW6N2Yz6HUT8ZcwZYPft7hP+aiA2WAupmyl5iQCJpL0X7P5gFKP6Pu1Fpy66G
ZpNzauwuaMSZKU28/IPNhnQuhfPxKFCeaP3wf2yPZoGD6gF6z/zShVYAfq9zTcswa2pNsMEH2EzL
RmbKUBMDWHeMoIOYTSiu910bfBKRgjKIx3oE7KN+Tjv/2E6f153wg4Fj16cPeI9z+NgwTTVdS+VQ
FoSVFlqCItsXPXdQQO6noCDZaYtkc085q/FNck8k9TJqgrOtbdwyVcQoUXZXcdFOl6qrcXGpZHWk
LCMF/wdTQBr+41cvS1+mJCon7FbIWndiawqhZgZybM0R/YC1hEXrqUUmobn4dPPmBcPUUeMIuDHF
lXqgUlmDWng1NuKHGs2Xzf5y+K8gLVXChACT07BGCPzLTY6XfQ5lgMuWVinCSrcVXV7Mt3gt/R0f
gYohU+bHqOtVvHexR4GHqOmRHWEhHS5SmcVCAOK6llv1R7VzWVO0jmKgrFM3w0XAVOTPgZ6VDehC
xohOOrmEui37NAzhhgC4nDH/GDAeOz8ySDPo3Dk/zJF1uUuTAaOZdGVLIRFcKatCTwrIjMQVr+oU
bZtVKCOYv8qiYFAVBQXSLaB2De380BSjRb4SB27uaD03aXszH/OBG+R5I+yc0dYc5rm50L/WnYyY
PANSUT8kZOo3I2EyOVcPOORSp1gTvJzmguOakjwoLwflvFABAwUvV/eKX2MVBHmSTTr1qPCdV+lF
lgkYVpYtbUSkEtVz/8vbPknYsjKIDml8LJGCZ3EQgu949QhgcZk5dDq89iB0dt0FJqjJbRT81zsr
M5Dh5KuOgU765jyez1/qA8GKxTxYSJkVBOmxt5Q7+ywgyDtDLlgLJgyiLgwxipH0wD64osAA2Cy3
LUXwlWLPwQRLMgl5cvXSIWZUTrX5c4s1K9XvSw2oWrWSiEzIPy0/BAYjsHGDnpupIftY2HFpK51b
Wm4FWBC+5EV4xOVx7kuyTPtBnUSckXhh0LKN+CGwfUTNCTnK90/Q2hEXdGu1VIk//CNESzY/Erl5
rjo6eZ+eFKihOCzm/LHHoxgONFCqGy7qX/NVFS26HwA5Xdwgx+Qwe6vlX7uYrgvusjBoEKWfpxkR
y3KlllJGiIvLUnJP8RDgL1MuefKd2nzQ6lUUp5q0H0PvB+aZiheTOV0Nfn8rnVpUtNzE62MyXX+p
7Jm3xrCaTZpXpzV2co3l9Lb+C3ZGNpo7CZY543H4BXDm5LRfl9EatMAwCoLWVI3IVMGi4d7ZsWOi
Yv49BNpwBY0uwXL4bCbY1s6FcXylRoakzytE+lUuqaWCdgg2RSnS07YH/HdopRAeQtHlov2U+wdB
wzWbURE93fUSj5bYY7p/7g4mFnZc+l5a4mVjVvmCRErB8W35fKt4UdYBbzVSafg59Z5OODKbqoFq
dAbcvvUwA1FQnDnjnuVHW/4z+WLbQCuUmiCuHd8kjbYiRIfsX3vYrZKOCH8evFf/PmeMO5Bahk3Q
u7ZpSbE+PUd8Jrmm8frCj8m5Zjw77avwLTTHGbLNh4NesW9TgaNlIZuRgqVc/6usqieMQXVT0108
tP4+Kogobt/0uJQPYzjoMsA1LeuLKxkmX47q14T6UWuL5iE1eEfGk0z0m4WS1RvWpQCLDg09cggW
lY9m2WUnBgnZMR0nVcYQVHqQ13cdtWREMt00efEqmOR2fW+zJGnMXX8DJBSmqhO4n+c5QQhUuhi3
Fq89XnxjtCgvcbJFxFD6YK5T5Ihrv3zOrPB6E7lG6dYgFXHQoOynmML06QQVCxhpYQS2eAq24XU+
VgvLezUi8zWGIIcyUHNNuX+BdvVzA0SvSYsnBmcncKxrgnWuEFtNVpvmJkBxpm+oYLgajXOaEEAH
DkbuEGoXVM/sodrFhqBWHaGcAJL1snwWe9Bb69cKIWhSDhDn416oIgaE5jZ36bWmoFmXVP6ooT48
KY98AducEQA24NTNJBqjmnCnH7iEkPHQzfxYIkw+gsne+wB8BDXMQwFYh2teVeCz7jmssfEKg43x
DyOYKOYCzaxYD7TLq3wb7yYJUkVoXCUwYMBt2UQOR45Xpbg/OZvkPgqrczqiJ28JDJOHYdwy64Mp
Ha2/LntXXB0Y7CUdxBs0fxjs4qkdi4Y3N3tVEKuAFNgxVFrkcBEldS0D4+niGWa4ujZYWkqs4ehr
dpFvtxbIZUgZKlDp40Xk/FhevRP3SzDMp1POv/ZLonVs0SxtKFGqM5nrHoqglmgLY9qUH4AghbnC
9YwIu5Gt+nwDwO7ZGHIboLU4h3mMHbiLHygM89ZfyFGN+5PuE8UxlJHMJdL+ehzGGP6arYKrzJbR
sU+8gd2Thr52JLzccpQpx4dzH2XcluumTuV1nUd3uAVYyHr6UY7v1vIx/qeaBCVBMicKoexnoRYK
SJLrGUaVd4ZV+78BS8Pk5RIT8pt6210UFxPOAJ0tfQfCtuGPFjHiuv6WNCJHKf19iN13VQmKpaiV
dY85a7X2IiColuMW10/77IIyy/D8a2OO6MEYj0GNxDKG79V8Hb3ZMW64uMV40ADPtwlrQ71mswI6
v4k78zQw9mRGkwSj3iLjUnygFr2N/ylcOspEjlHuLf6lf2asJhYiMZMdfS8OrQj8HIAWC3hSsnMa
tzDhZu6/dc7qB9h6EURMwQ58Sa9ONYPhVV9RSlJhEAtchXr+GrrSqLutTsa0mSIOM6XlYK7rdCic
Lp13ZL0KyBpIh3ufWc+yZlEJCL3dJNAdgm4xzPZwpymOh/Ujm5iFgS1iXrxcY/STA1BeFguaJ8vI
qIZehqO9sIqetrcHHsl/DO8S49G2GtlUzODqk5yBp7eVYSPPFKy1jSJyxEoapUQi2SaHepL9ghAY
6DL7+MIU3pty0kvXccEqdMaOT6F93+HfwFxxP4N3ibc8KuImiVAV49JqO+B9WIl3UOg8OVj1RyP4
fkIxMgvGa0nnzZUXt/tKzndfx0ZzRddZGG2BYbK037GKmAm8mR7gOUKgLN2HjXgWdNUF2O4ml/zy
I2qIZ3SoNo8gm7/Ha5pxdALLL8zcxIAyUyviYLekMCvul98p3mxP6EBJf85QNBOZqa4uyGxWYQpJ
5gFEqKQrApGBE4AQ8bmZZyUP1qc7l+lOcKOIiN24ydG1qeFfYYAddywMRhOw/2Tot26KVtDqsL6z
B2MxTY0ESoJs+DG+XibmprIw4zWomvgEXuWr9naDkdesj6jd2gmrWa+gassZf5sfVyNjutkIe8GB
1vFMTWxTd/9rKKAtP8THviRMItIUQyItOh0DICKkKNYFshAXs+iAHFrVaCXIXy4iFqoG028bBaFb
13LK3R3zeG22l+5oOU56PJv1frO7LwvjSReVd9vVEa04E05fnZ8/IutaFScrLkLoSqv9jYMQliV8
aCO/SDX3rLrYIFlUep1mXTGD/K2qKBn2+1kj46ReYSAhzMij6j7e0jr9J0/Y7gsnvIdAE1tnS5bJ
lrME554xLX4QDhl7Vce/a4atDg+jXkg9lwb4uu8bmo//iXQrSvQ5R1N+SNxvQ+/ukzB2knKq/P5y
o/boJbS+padDgF/xTCFaNIT0QqbbtHjcilYHdW9hbjsf3xAKEGt+PKNyycFwxasKsF6rTEttIjnY
e6KPRdZqZ2tiyUI01TzG2qmYZWqjmgofOpan9c22AqYKkT/yvU6D4oMJ/gJ0z1wpJL/py/KVjDci
5ZtVZjKseFqYxrqPoQaZ5DpwpCMivc300OCWZx9CvLbcEJXsshilymMfucP2/3P63AESUP9AcXkg
l4PtbGVWP93XpcAqhFdO/GOj7MtlCMReRXzbdGC6PrmhSVy19tvQ7zcNzxF8Xl4mM2s6NE/UFaQc
huiiPKIs+Wb0/H3t9cfVbrR96h80CUc4RznO63VZGjQSc7LlkpW4WyeWbhfSl+pp0/E4kt34iv8x
h5Own5dYkJdAf9dORMUnrNtSMlqqauRBz0oGwFCihQXbsV/AHUdt58oCk7PgOZoeZks1jQ52aiSv
18NVd9pWN1SKDlZDV/CcCZ9VrKg70DHx1R4+8Wmo098bs38Yvl8oOwYV3vPBLaWT/OffF6qjqnlW
jnRcY9F/eb0MiMzlT0ICx+T3W/vlSvc9hjKNKRRRwkN0ET92Z7zPuRlw2vqirJFRktwxmVt5vTPo
Skp2flSiROMzIiiDG8VZJ5G4wT4d7pl4f5EtW9CBAEpP8/Gk6/FTLYc56oN+76gQOUzhbpr9WNTb
DFclBAsMqNwE5s5sUmXaAOsGOS9HYIidF0tpGezhjf9RUYtXjqWSp6aokpBv8b3GngNpAg9oKfRh
s79eRZHNazMq4lir0oy7ED6V7jeIwl1KfPjPx6IJl/KBEqDsgcBkMZs63huHIcgrKhHYQBmyfNKA
al1lbodeTw1nAeTWKBMkr407/7OnR/KCy1U0kwN0p4g9EUrmPmA/SuRzptq4k908uvR5BGmBLEsn
TxPO/WyyJswSUh3S0rQAg5VfhAm3jrh9tt78AGcALEfgXyjfhRJSxhNpbB9YZ+pXAmoC96B+fiI2
mbraPQ06jynMDk6sNR1fwh+k6550rmXPTBIK4VAMclzapzEd3/F0GlRWDVjS/7j+kiyl1i7z98kO
L1x1rqt4L1ZjMrWJ2TcjlGs6jxuTA6UtVht6egyrBxPqM12eCmNvUSTNO6eOS+RB7BtpBLJag1dh
WSr6+iqz+42aoVyAaADxCHEaxTdkVGj6V9eJs2GRAxF89bchNj8sppvZkOBhZ2hcgG/AlU2/yZH3
GmhHAYClVjzU0jMQgfJT3f8asWWtkzgWzpFprMBRBQ0SFwShL4Doo7BOwnCe24EY2IRJ/cd80fCI
nVMiKuCAVfQlXCP9eIIE33dXhlmTA4q3/AANK+FyQ5z2zNEcO2aDn9T6phPJZ86a+eDU+7khJqnK
Y+p4z7uxgOruLBcti0C0tzICpNL9I2GFapx/aofHmKHG2vMr7k50MsnkyQpktpTaHwqrAE1xVph1
SmVEV2R+9dgaxKBP3xGDbXHTt9ICxtiLqQTmcTqKKEM6MTNiOXe3kcbJIEdV6yM2FXBGbvBV3VqS
E+OWvDJ9PU5YIgbRRhJXqIN138ro7LP0/QMUnsRxoxJwTxO/chdPchNgqRgH5CUj+ZfOTNlU7GFQ
cP/PDboKd8d9UFnCwanIT23serjBeyJCjnlVG0STNbnE/f03N7VY9cq+AhGlG3wUEHdfy1EYgugJ
e/z5sBgDcx2x+4iaXGc8zy2gOO52i/CeYO18so9A/LmXFtB0R8is2AfWBrBXrLCFYcqrtRowUh0l
d/OTkjsWqRavZbCDNF2b3H8i9nHwmNWzU7uFHfk8UOzP+r8Yeaj9dvOvct24bq/nM1cJeNhcN1oN
iYVN5JdEAk9Ix1TG9tJEp9E3mYguIQMTy7U75WaOCa7fQzXskx+e+9Raet05DFmXm/Uhh9jl1lMR
x89k9CzzTkK7dWfcVUlEc7r77DBGgosnRF8Bc6fg6Mav6iFkOOBi8j+fPU8IEDP0PL6YvUDb0Kc3
1ZaeCKCmie7oQAvfXb3PRXyAYXC6R1CFaq94S68UbA50WvDdyTjljUDrygJKIlxIruDsr04QpzzV
viGKEz9X6PgXXxtuH4p9tqMhFtRiNW95Um8amcna6y20jGhFzP7wcde8Ca8Yx78SZSK0SurHbgR1
OFE8ijLI5jMo98vcDy5xsRCrdYUG9G3Cc+wzQXGrCoHmi+johIO3uk1QhDGf6PUml01JBINrRIDe
h6o7Sk7dUu5sARYf55OK7XaoODzW7YfDhdgnmfbbXnZlOPZtHUGC2VQvnGe4RMpzqpbE0fIZ850l
tPS/ffZTCzs52tQCsz5+Y1v1cq2ME0qvAAgb0Mhy0Pv11trH8OkoZuGnoaRTBj5wD32y3VXYolEp
Vti2UtceUpLJ3zzSKuE8Llzw1c6fPOkC3ziGtcG5zUZdmuiXsgCtRf0ivTFnpUq57mfqfmfkINEH
+8JvZUc6+CXoxylmzLiSq3u0uCrOrHB5tI45FK4dLu83PZQnqiBHQCfsq6Xq/bsKBSYvzU5mnZo6
XQHhpPzBGpCPspmivzcu6MJgxT16IksqGYdutzWMnBOBo8MswYnN/JK8od0AHzZhFx7YlYRookpp
EAt+qy/P1bmTOoYtoO5o+xHDS+N15nZAGJv/MUQS6ed4nrFoc04Gfd/yy9P8MoRYtJkLzUY3xTuy
zF/4ERmnRMMxH4C2uFFrXxLjuOhfw8nfyrxuEu4+1+kvLmTwiTxgx+xbi8M1yRw6ov3t62DH9KRW
Z0dBt/GeVaZOGFVj7STNNAnBQyC6x7zv8ClOPMtg97Zu8MZe8UhYdMWF7K9oNFZ9FLsQEuDTx7ur
sD1O+eeNBFfiHv8Zg1VjJaqYa9ylLuuMt5MAKW6jYUYfs7D05iGLW1+Eih46virN6n3eFRRmEJLS
FiGiXtWTKFQjhCHHi9NAlC/Iqb82ijXb/A1tgY713nm5snBWbEfrhaRxEWEyXUDMsie/Xxh0SlX7
Ho0DeXfAinqaz6Pj4kBb1jTwTtw358aLww764wbf0qVa65xlIsNf8YwaSWiGskFOpJNVhmPkx8Ye
cH1yjc8cXmQ4h5oz/BMnhenmKFJrAvTaYTuUO5RKL41iAKTovO8d8cAZl1F4vRVYSu48mqaiUOEq
j9UgCbHTS2v5qJxx1oHL5sJ452iNRg7E9J/moPnZg9G9RqWvrTsYM4e0XkldEpd6BbUv8YPsDoTs
FRaHtPbbGclrrj/uex/OCEnGwAlYcMAkTxau3HjeoVD105YTXgUJnTgRsL9nztLF3a8B5HMhodL1
fj008IQkiQ2AXw7hHzUncMBCM1h0Y/RBaEn8vRZE89k4AyopRPFMp9dZfXj+8d2v60VChcsK+LF2
L9CJjqPlP/vCO/F3gK6OqNJRDpQL7yH+nWPOzi1JEDUgL3sxmyDU04bb62+IVQAxjn9nq/fdjjew
HjUl1XVkUO+ViengS4tWOMqaEwFnewF6tLSWHmbBjLgKP9IAFfVmvqBjWyFvpbZe8cti9fWrdYgj
m2R53BUNsBOe9rTduf9/V0IQN6DrCfd9zRTJYeGCyf7uj9+hTphmkn6aNBBF19o2B2r7o47ZLR+V
Izkox8WvYDTE0z/F74v/YTSlKgvrhFAYFlQItWHh3y0MfgkKfrv6Z6qSHAHbJ2RpFZElPhURfWTM
4Fy1t01q78QJrpHnJubjqHgs2rdtU7ogwye1lBJjop1gxp/NQzsX1vfbhg4lcENqRhJASQ0BKz/A
DgiTJUZRqIVfxHphVFMU4G88D5wzAX1UdqmMg1oGlK9WlVq8uHlRvhcxZrYjciukfCqcmnZlLmxU
VhfcawfswXhPpiM36w+TBI9AWsvGkHPUqvErlNOGVRY4dvzkYH4QJf6eeUjlQuB3GqexZTzxb7Q1
PjhlRsxifzXOeipMbVeUIbrmTkcx0TxZPFPN0mI5KXAyBINVGGWLhEg8e9tL8+y5gntLCWshmi2V
q6xk0NkCrY6e44AfAGPBHl2E3FTXuHIa6V3FqpDjqI2b5EFPQ8oCDro+Fl1kkV1DGU5/IWi/bsQd
BR6FJ4eafv8NjOb9y6+IRMeFmeKxO35tEttBEzq2o86XCBt0TAzI2ru3SK/fg/osOPoj92QqL0iq
t3TPQuZ1guGevfKjofBmJmybSub8OOivAiZuy4+5ZstECCkPQ7lY4nIHsTINAIaWezfVBjah8SFy
nAA2kMYvAwY4RVZy0JaaCYag9GLmWcC18CiPFHXwv+9kBMFwwHpkuskrbn6lqCCs58cJR7Xzxuyp
NVZP8P68T6YUoM2JbZLu1CopOGem07vjrcXamS9B20znEQKzFK0Rg/J1ILe3TorqAvkAnyzy+xLN
nczz4nMiPOErhHB5I3xd0+VC0h0mimlJR9Y4gVOmWkJPDyV6VtuyQ2IfYWsD67n+g3gMvz3/cb8C
wBBrc5N0LB+E5xx74KeG47ExhXg1DVL0uuv4q8163Uk8KUipxvAXrCotafA8/kxKA6IFwpMMgxfA
ULmLzc3qcGxkWW5Hwprm5HNEFhvjUBFnNhqtsDBQUmqaTV9VNs6/qnAVTUNmJ++HQFzoOyq9mdm+
BhVMdnuDbo1a/huqBNZWdoxe8eZ8XNmZ1aoCUlTIIF2mBsh3Z5T3g7Ud/8saKfIesspj+FZKcXLe
NswU6NpweJGUVtFnOlRBc43189/f8Bj8G5eH5LAwPnnDihPngUkOGNQ6QXDXDJQjo9kAXbhxB4IA
Atjk3uVNxddnkxPs7n7iMZuRRu0xAKjjQ9k6WPmHdiVLjxkFrYFhTgMCPtS9G/aZDtwRkzxlIiOw
a1U8bnv9ZTyHqnOeDZ2QT9MRtzmHIj26PNVhdGxtyOJ9LKNgo1hvKQur9G8Yl9Rb5otlDrcFZDUx
VB2uiG1Y0C3OqESTnmgQXRUXow4jtMquETvrR7soo+mRzcOv0ssV5OpePcKJtbqw2ux5ipWhnHFP
utX8njaSnsOmwMlzJNLH49qKxTXt4BfAGAZajUSDvBxXAQOGOnjQwnDntdBNdRL4ld3h2CML1BnN
ivsodKOo+7aSf7/gQe/99s4/1sLET/PwV1ink3DcGlmQ/CftXt701/k7LrCGU4Hj/AVM4elzmk/I
MRcIjce9IFIuxuWjS/FU/w92/78wKawBQmaFK8YG60EjKO3GDFUXjB+CzCkhAhRVA59Mir58dhHX
WRlwX++fCXVOeaPRKvwJtTdLns0XdLfGxif7m00ag6CuDxJBatV5weL+fVxFpnbcoWtj/0BL+sAo
tJHASvogNN8TivsoLpdAD7NiFM/PfTbVOTRcXI96a7bK3Aftl7vpurndNyqjK69rnlsfBPIjgqEi
V44UvVpdS/LBOtgx5/tG26pJ6rL25gjgQqyJUkTj79ttBqCwfcwqjtThGDsNunkfzG4v63+BQToa
Mr6SM+8vYNsGt28wwda/3ebDy1dBwEnNQpWrH4AFIDkSM/XEN73IjCutAHygVb2koZzcnNNDlIlD
pwdyMMvWBdmzedKK6MizY6rdm9wdiXWCGOQ6t16nSCHnGa4QoCSymf7vOs1mKUytxcgouTFlcUbc
9o/8+QFstmj8WhQzVmFs7luqQgeu55Rbuk/65I51xg83cpYThi9boRS8cJG37mCu0boABp/iGtsJ
4l2RQVmFiUubIxIXNOdQyaduC63KhosbVYiJWNUm/6Wgq1wno0qSubzrSb+Vq6/fpf6Yj7JjKxnv
WC0KrWTbS3t6eKI0DkZONBhu9c0uA9n9xEbJJ69aUxNn9oMyP/KWuYsPgE2oVj9MWOCeKncpz+TN
fwJ4+SmBH0nSMeBsYm24bA+3E35d2DZpFDkfITYIXo7z0fDQhqhZz/Z9XVA9uQpD/hmyxgo88yFK
e6rK2lTJPrYSHUQkz0phQzgItZBb59iyZoDRo3T6zEgLEyiuM4flTPD8nig1jptF2nmgEHUXL2F8
/rkrizGPXqkffks60rl9OjJAweULDMdnqXuOZovKsjRujqBnoC0fkyBsRf3bXjIS/ex9IxHwPoIX
01PrxXd/LV6HEt06d8Kg+NDPjVBUTXizMoJhBfDqwKyEgjF/BFDnhPcHzVai1b0388T98uawe1BD
K0dEDFCLIWypSd9sy0YHAy5gorDGrizACR9OKvRyZm0nsIX+DidGIX0J+KRbByi/aW0cx5eV0Mts
AoE9KBjanhWE8wNcUcwtr8ERdwriUbNSMOlpS/QXFIQoBvcCVNCRw1ItHZUeTlw90CMnhYm8z8p/
xFe1r7/Wxl07ubKLSZ/OCG6FkiXMoC3JLzBjX+mGFSFHHZx2OaD1kT6p+ToSEZhPczBfSH4TqoO6
pwefz0bNJMlGeuBMo/dNRFHi0D21nERxeBLdyCMgabMkMkn3e5GVldtVlls9PmK87WO9YgmUmamC
J6fxROPht64g/7TBgVhMfcZ/ViMBXtHvFILZTDU6mDmRYjz3vQa9hpBLNiSvmKxYomZiIGrhFHM6
DkimyXn4DY4jcQ6kmkx6Si2Pkf9lFEY2Oaji0xFJIr0uakIUuleLmCyMVFNQhyG7Hil16FMJh7bB
tdFR4FQAcxh0KnMVeu2i4NiULkUuRDypdwE3ibZMIr7vTr07wAoz4UOLnyW2k6afp9+EusdUes2L
643OjiUMG2QUWeyVkB4PPjZI+qLX9eXQTvLvBva3ERZVtZ6LnGU+TB9/mh2s08bnNNlzpqleToTE
uEFaaCktkLAWXlqJGaXiT3bd8doFw8rwQgwzGAt5Nq1mg3ayBZbxX3wHKKFNtjBg8CEIw7O+VlW6
Q/AYrnthOKEB5NXvdcjLc31t9ipB41o0zuWrWup6uP6+k9YClIvmrWcZBKv1z/bK22DvoeQHq3hH
wX2KXSIIaW2EOYzeET//42cdERndmcJJDPXjHsH1nMoXrjhJrpA5OfykF9x79x/nS9gvQ2M7HdgS
w4Fneariuuw3ljhUL3MdF79ULYKIuF7DroYYuWmrAV9H8ONoG3sPhXoZ9K52KI8nVRc14UEBg2ow
lyHduBGau3eIitUeHU7qwVV1IyGx48eR1JsPqjivtwOshV+MUgZ8kFSBs3QT4s8oWny/TglHOi9V
SXZCCj27hZV3zSEphKkhMu01DhK8M6kYuyR4TFSgOUQH5IWCbAt7xLn6Alf53e1tubeZqdEklYEb
bLaEI1CuJCrBMqzpCnqwkwhIZYqlCMik5O3aRfzztNR48quin1aLxWSTM9vgHdVO3KFMf8g/gc7U
nEH+BrqDuuxt1Duconk7HZo9A0YFthdyYD2Aa+Z+kZLCG+crYiKFmzJUnXoh+MR7iezXnqc4KlRK
GWrS6xn10HSB4dnhWi4SkZDjsljqQf4xLE00BfhoRopzTugS1a91mj6uiOel62DXLUXlbmFJm3n4
J2FPRTOwCcvHipLqeXuRTHx70dWVcmYfzvlvEMKtvB1uccuW0HSAGNaFE9DHcCg5OGi+JkwLRdkp
Z7TwXBEaJv3BQfe6fm9eyY7Sps8rxOMe8XX5eOT6RCC1+Gwet5j+dOxbBPk+075C2lRCflvit/1Z
U+XUtHPnzj7d5+z1YIg+zCg5mQFORX2lyeP4CXpPd8s6Xtk2J2VYtVygRUBf1b9N9hpstSvLN4uU
u+F/YXnv522693dgaU0PQRx+/lltHrGbaPp+Q2VtJrlFMoIs/BZ0j8zZofkzrO4OQ61+QVq4ZzHu
I6vMTCYBBsH2i6jiTdH81jr1qeG6cmLiPZq2yF5sYoZ4LDcus2eGf0OwWG5F/Y4ub6WkpaSREgF3
eltULEh7lO5hgO0adiLJyE8l5W8XXcVXXz8JkXHOqEj21XizzwvP/wiCazsOqx74qI0ucTNQ/dMI
1BgYOpjqD5FZh4SMmcTotiHW1pgsds0SaWLuKMlKrx8lofCiK52OtpvWOPV4A1kOFBlhUiQrIIX/
WbeOfSJOOaqpckTqwCkx4DjTZvGqP+8MbXlONwcZM++h3j3dMnnZoFmD46A73dbL64OK7cG9v3YO
8+72m754n7I5J+3gzNBfeM1udUyFu6w0WM0tCfOEuej3b9Ya/4ULJ0UKmCMdmCeZSosQFi+6aqpm
4kYaCYDNtBR3yuYXcPDVrQuAgpvGjvhEA29JoTIOTXOHu/feL9DWTYlNwu9MkhWWYljwGDS6hq4V
l0W3/u11EQNRHlwYmEZZD8nOKASJ5ZI/he6HSOXMKMJqkgOboKR5RHf+nKW3VmH5x12XaPZeaaqn
DAGHcFNyRazZAs/Jizak2MWozwX9ts6orS/qkfDH71t173jp1lN1tC859/LnTrXpfM2ALORXvXhM
uxviJuReimxhD+dLxXVcqVePQaKsYmHsn3vZsv1eTLbfZi1T3t9+CN/RFn+jY1d7fC8F/+XuaGGp
h0T+eyn/uMgPDlPRKkb4oCKnDs0Hkk1/ThkrxKsc8tiyaqtkMnikMqcmaQN2yhGl0npVi7s/U/qo
mdDK/fie5TOWQle14MOXRVi5q2/kkIj8m4NQlqnyNtMC3jv623tXdqZmvcT17jWnN4C6RdORL4fs
3aWc/ipFf9Gvw8NIGLN3IIQ5fm0tUTh0sOx6KtexGmrShl2XBEs2CUHORovBlkBbxPiwSK0Zmojt
YURe1gCZt+c3kZFL+cyOzij7EWJdwjuB/hkEbWMfVwRDb7mCwcmt3sUWzCQx5M/5ka6Cn4AGtAEz
0gVfuyzFW6/BIZZk8hNvBf1N7IGQ7LJgqvUTpU6b9LMOHyqDX3+66Vr00seWR36LObny+9Rg257m
zjWzjsxEx/OB2wwpNDRArWThSMuSsn1sRlKP7mySEQyskr8bx15+cflyU4deMFmxKmZ2FZQOD6u2
AUGl07iqho0YvLsd3LpRBfduDfrQ+YKkjk2aGnjHujnclTMr8l6rFceZklve88w+XqaKquJtVuzf
kyh4Q6Uvstd4DdvG585mg5g3aW7sXATBb0rThEtxQ5P0Qrz8cJSSBxirw7CZ4GK31q4g5auYnhPZ
29Md/TwxxYjPRizdeKbV6BPdbggPXqvKg9+KgcQ8UQtkDyu3FbMhH8t0zCQ6BCpnuR3AsBMpbpDI
hiJ3H4Ccs7GRRjTkd5AKar/r8Cx58ixMJ41uen4Katd7H9Ibq1gnlymOolGN6msHq4ukp0u5U5RS
rPRQuKbKLpadae/qa1F1+nL48jBw33tRwoKRLpZ5zqHXZQ7n6aw633xrf8LbP7xoTy9Y0Ts13hZZ
MAwB3708/b9dEOukScAie8IYTLVY2hIKHmAfEEIgmi8uG4cAZNtO6MiFJ0+Vzu49+86fJZLEMdgJ
6tUn8niwN4OrVlNaRdhwRqijRXmxaejyR6hx/RxtaiQAA8hto1gmfrMPRuHJhKs71WRrB6EgnwMB
+1DQYb2h65m2A1WnHgxRX7R5M8I0TM2j8ed9vcao/Tzy1ubsQRhS+5BEjKaKR/n5huhC2GJPAwhR
e6xqg1qRLB/xZZRj4gdHsgyIYSYe5ty9b6kul2wnOM+bhS6w3PDZKRFMD3x+HkKaNk+7OxCKKcza
BUTSwZ89GmaEK0NT5u9M19vSceXnusPNOW3VzkQ8RnM+65dgufto9Hx5uxWuhigHxHx6pOc9lDy0
VPFvwaRgBRXV/AlKuALSDGh0yVxetUQiNH3XOg2RJZSV2RCPNiyWPapkv9h3ohNUldw0OLlSJiBE
JykkzdflHcA5i5cl+d+3jRKTMRARvxN/Hty+IYJcr0oyxWic9cOJk6yWKsBxPx9fLfls3B6OoIbC
g6QSkWhRompak9cgRUjbntqTCPXl4qTy0IcB5gGcCbGfQFzjdgTEozkO+KKrr4YeCX6IgiXAMdWQ
+ZPGc7+jbs7siUbclO32e3xDTRJbZjTroZJHwXvj+aiZ02cCd8Hl+O6CJAagy9ADuxRK/IpIpGUE
ZB7qX7KZ0ERiwvOSHWCmKBxg3c65EcPQJEOMMwhIwlgUjvc0uwMc6uiqY60cPFYPJnunN3mqX1al
s89DVSF+qMtyhwyybXg1GPTfT6CcwIouIbTN5UX8leuN2T4zlfNtFusGfnTJBVJUqjEyWYVthSHB
ldRgxmPHZANGUP0CnYMFIgeR+nkagXZYP2Qy8ZZp/zH9JQyteIIpS/FVNKPnbAyO5kZRC9xmcadZ
P9a4ETJt/CiwUp/FejrL+Ypq7gGz7AGNNGj3sQ4RB6toVTj9Nh87v2g93m9ogjPSGAC1rcDBTeCO
cfbVj7GN9frvIGQ+9t9TkqmcV/KwnD1VUN/c3BYdQsaddtSJ5H94lFbDtTHPtJ3cvvQdp8SWfMjL
oLGeZNDmOviZRyR5SznJzqMG4h5Onrsij1XmZu9r5nEa6sd5YMXvAthu8tYNSLgW2+h+4dg0Vwl+
rpmK99Nc7y0PRIwpi4tMH4/NmuQXJ+s24aPz9x59su+0iTP508AtrwGwLALff0fUxzP/6ZVtE/y6
w+VRmlXdDdtQ9J4dIAIY5onddiNZwKMIoJRInL3kEhPm4pvBsgjNE1lQZbC3SKuG9RQ2A07M/jHs
nKIR+inU8qUC0b4st3caiIf1QugLm45ni/IlwMLWy2Mm5ZmR/8oHfFuCfi5omyHAS203Vr+N7S2h
8YPVDE1g9P5T6OPgMHh/X3XUSsEostr7ajl/Z5XHHwEnbMww9XFwURRvh8PFDnNVPGSo9H1hJumr
pMWfLBZy5EU6BVI89aO2WDbn5IjeU+iv7YNwFjxqoW43uaNFuG5sk7XgWQg0A1U4ctG2FznM1zKV
udcg0zpLJKecx/PVrQ8tEvJmbsmh5OFbUMDhuA0B2HHsFpg2D/mkV/KyhpSKJx622tSoYnVOTmw5
PhZ9279Ux5/meAQRVBGbMuzNFrWmp3AX3HF0Q8e/bFHbn13mBBTqh4RJHBv6eJ9XEfZzOQqwpG/9
tIfDS0ClCRznCx3v9h/sTp6EIj4jl5DwmlLtJyO2smxep6EPDIOoMvXZtkLddeppCRToa1M9p9Zt
1fnjY2wFXdu2T6TeQT6QAPB2elgMzr68UZL2ScGt3RgIXzaq6cUUbdx2EEXieaJ5CFsAZA/AfYVA
suFnUAGqlUtA7Gux5aaKLacSs3dC3vMjuzzcJDb0vFuTCoqbUFNSZA7OiWSZqxf5CRm3xqepdQZQ
awUR+FPOBzfkCYuB/k1lwzOY51vwIazEM9cbnvAr/P1A+pO2XQGkg2TalU4Y6PArT3mkceZsr10v
xMwY/UTe0ZjBqfPfenT1nPwIh9OvfiPfzIv3BcKzdkcGSeyjSXuXAI+VlBNgRvaXhdMtBl0var3R
7jO11VMOkIGlNiQgyv1e46ltqJ4PQhRj9p68MCUs0xnOcBQ8TYpI8MAIdIVS0DyKB8LgLTof3Lvv
WUrokhiZFsPUevhuh2JqSPKsP+FHILZkFppunfZu9zzPmTTbHoQAuo4eDXV+S0IkC6TFC5UjOROK
TMz9trUeHpW2utzRgYimceSU6/NPvx7zSyHXJlvRQO6K/qPYRxaV8xr4/jbcOViciOWu4YiqVbDy
o3StNXNRFAY2xC/HXo8qoL7E1/BGYrc/Tv5X8ijR6xXeEK+MBd2OXYLAkCNOzbO0oe0gaFTniQR8
UJpy85HvcrEsaiziMiMgIn1Epy8pDJYh8fkYClECCKdnw+PTwvQqaeKvVvfRLeCT3UBz2dkTGaGN
CgFcbeVyH4rRCG6vTug0vaKc8Vpnml0UHqZfjXfvFdhmOUgNCVX1DnF8uYaHSUkRKckJpbLTFJz7
DyuVQeNZuwLhmKesha7PpRHCEaRrdDfsSCVcf1f5TfGxAKPDFwtkjf0zaEVBsrPfhzKGHdWsjIDM
dqKj4W5woyoqB+suMaCDu++no+/qNtoDOBZ7wQ1RZZ8nGQVQvF9YRVA8q4gcGdM5S0yYcALBqcjw
TeMoLfuyFJyQrbAzi7FxMoULEnnyhMmt0I/nEulW9PnIZEQuv35vTFoLH5JDt1zvjRekvZWyHDAL
jhQd9pudTE5NmZaGLoHVszoMpa+V+eWu7eD2/O6rm7Xlt6siRrtAeekKrNxfW/QDRRg1T8Qzty3T
yijqoiKNruFLUUWDrctAzzeyVNx75K8btVoKHJwJXmln9n+I01D4qv8mL6V9X4+sYtQg0iyowiVE
MGo5wPuPrC6LhRl8CK9/4SQiRCIfseSXGGMsPEylWbpIBcyB7MX4+Qf8ALue6LRfzmGZLMbONgab
kPbCTRxxiksusgHpF3qd2q1q7D0tdS3FupPos1UuTEBOpcc5sONOFyztlO8WQSVOxlf18vO/GgFl
STIV3sUNZ6V1oRlkA0Vscn9BdqVMtJrDoUJ1RODncIBSAXOV7zXudI79MEIJNx4KTqnmva/Ze03G
S0fRot0OCwISjJ5eQKEqki9ClrOYDbtZQ1PjglB1EiUvQT+MYABDF9xZ1aTPDUNgYLAF7JecVJ5o
sW7BHy7gIgsKcw2kNi8+EGKD1QdDND273Zh4j2VP24F7aJ/AKcV+KGQa2+Lq8I6rc7mL6Kbbl/er
GMLnlVccVKB8xnEg+47Wme1GTiHagCp5umbw+qgmtwb7OPT3iGTZOtEiS6tw/ejfxg8fmNbavwBN
uGyMxAG0DIvpaZF/cGy/oJgCCLjbJuC9AWxVWx2X7clx9ag3DpSdHHl7dzsuRGu981/h/KxRHnVg
NpLKCmubD8BKFkF8XS/aM+U4Z50TTYGsSOHTXqbwhj6ZTlgtY36k8J/TUdbk7QCHS6/72+Syy65n
HwXY8xBKqyfQsWHffU5WmWY1gcb57IPZtRfQm/NsyTZ9YjNCfdkVm/wiaBQYlF3UZ0VOGpqarM86
+AWhhBQVPpERaOlBKgOidNXQktXtD9jFPsU8He2v4nEi3gxrNhJ6nDgVZlV0PKVF16YnQ0El4dh0
YuEnniFxpjlH1OvhGPemDGb5nN6m7Fp8wnbb4Nl3C9zA0P5mwZ52ZNz/NJOmVWjRb2cEDUGA3ZgS
v5/CfyQN168B1VcDSuKuKjtUpa7mWMxa0sYKlEQojPDIbDQ5sraBhMoS3MQ8QFRxCavE9iTeX9+B
nDlCc4RzUDhm2CnpWC2fDdB0r7UAGEDfgsukU3Gh6M4HA1/848MWtfMbqYeAHplnwGvCneCBOqbw
0dBnmyz4Gem08QYyblMkq/OtJI/xur/zjthIQ06s0IJRi9ba/KkOwJX6u4tO/vMcN3UN5C71ywD2
RxkLBb4wWD7ZiWpGXeR/jtTG+slnB8+eElnFctcA3xWBahTAtRP+WxCyXVm+WyLR768v/MnnFmxl
pV3gSf9cdcZUKSobtw2je9JrfVq0jq+TWlSYXQxyFavzOw7CwVQ5RzNjYs0Ck83exs4NnkWeHxlm
15XVrHafVD+0SESzUHG4qtEYzcpK4FrDO6o6gSAzstxhahKDxHHfynETDBp2rL/8YO5OEQnTLlZ5
kt7sMuq258SVyM4dP5tYEZUolfXWCU2do/BgcCCoJmTvh7OrVCBSGmNaVliW2zad5e5mmZuv3m7v
G4LU20FP9wtszwVGMXdWTRwvzjyv+CjqTmCEAYaG/3piidRyTZmgS01fiN1q4mED8A+R74zTaAqj
4LpQCII4LiX3mLHLy+P+R/1GCpYX0m4AKf4BlQ9HU+l2Du6OGVbVnc2zpwjiy8/bf1O2B82BnFJ4
69fkONW8M/J80zUOaPixNpo2WThuoCp8x4Ul4hgNVhbGcsMzGCuqjs5wSnk46xZz0TxeWI35nsh5
n+sYhOzLLDc7oW2T5zvgDF3RmGYi//vAPVbofXI65HOR44ZMcXdRyq2+j9Wkvay50Y9ZrWhvfmIN
kXrT2vQdZczbIxK3MRvTOi1TZorPnWQcm8WCacokPkzZLDHSUXG9O2dOLAKUqWt9fwR9/yQJIg6t
m/+zQE0sDy8uiQil/WnzLqpTU8yBkMJeTdFHU1Rh2Q5RrK7O9FNBcBF3U8NgMYdU4Vgz1iqzcZAT
T5COPKSHNE0bAFv1xRpe8Qh5wdYZ6es6ZnoN4IARDY7HL1kkAwnJBXajyfXWS+DfexSL2x8GJKhs
VkgBDRNR3O2rOnn5slits2N9WEGvBHoK2lriauku0wW2PbrafVAxKuQXqYBaiF4NN+Ji78KZDyRi
HIDOGlL3YAN2UEkmjZ2d6dVoQJTw2a/HVqgAh/vCnGLaoEsjcf4Kg3YqqCCvloEDTLCcJ4hm1Ibg
lId4VUavT3UhhjHNsllZJbeayEHWdro2MJaKSGDG3dC0H82wnRB/o9AHJwTN0+mceRcUDZfIcnmM
29SVweAv3AS3JOpAdFnUentcOqO9O+mznislpCB7iEgidggXtzBp3WA8nL+keuU2SRXrKlywFuYk
s33PAfHfMOixP0U6RnXnzombntgqUanym68KP1qsJfnDHK0RM5mTnM/Wb13weT42i/u0dMG5zbGa
a9OcLulpyMi+YULjrOJ3xEMc+vD0jDdGO9FgO/vJj8T0KmAyPN3Xnto5rBMwXQazGjXBDD4WgHTy
A/exS1UKXJNecJejGrBsxMxMZe0Pu2oKkJnH3/yD73ojlzoJRLmia/x8TPyxaYAXA9vyp+M73lCy
kJf0BdSTgiRDDSMFIFOFkEVkg94uu+ejtcxP84AferZIbLHidTm2r9y6VGlqS8i8BLHsm2VgFPpZ
p46xY6Wrw2zDHER5nmv7C0pHHntvMAQrsxK4EafvVsSdjHk2HeIPESGaGLcdy6nuQXSq6jYQITcd
eKLLtdUJtlOxHSldjh/8m8J6ojXGIBjXGfxrCy3baazZkWg2qquLdyNnEFxU8RjZwQBTBaLeqsdq
xJ7Gff5Sw3wv0gWS91jmJ3ovw8Im354TJVOPVDxjfRP7Cmk702R23xVU11wltZD0XWMhFFLc+Iip
J6KW2b+l0S5IpfYs4BKTkWNESzpJMTnSKyAUK4ZStrZs+6d8pkR2v4bQdke/Cg8SXAsypriIwbbT
MfrMt36ivRjoiSifFVmQMLWPcps0BjDfjAcJiCuGEi9FoGfJwQdEvQmbRTF1kahpfESdFxDdVJn6
kyQdxe+iAOqwuLurkFrVUL1jKapuCAVnBG+tCy2yMUGy26kaddVFim0gFbQZuAndI6y/Vz9tF8UD
vup2upoiJhoj6uukeHSh3mX7x2ajunW/PHtnVq5FVSd6cq8mCpdu4dCl56nj2RlpC6LOxmeIl9NG
troIb7IQ5lRIbjNwjsmyPFIfyVh/HB+HeL7nOjm6tb1s0aagSObNc47jeIVwaP0kolcDaH+bAOIO
cGQzDpQBqYHG/H5bzh896irU4Km4IOqIGJxBTvm63r4LisTjncpCuQfNtmuB93tHJhuB/+K2ymfW
lx8WL/gXCZMVi9urz3Mys940v4ms11nPidPj8El+JM4S9PlP/afvQgznwyh7GGW8E7NWtoVbjJ9U
ZvEaNuWpzVK+3B5M0jfCo5DrtQJX9fDsEY6CTnpMvX79nnnQqpRblLb9luy7d4hEQZGFHK+d0EsI
IoUIHFIf5gof0plAnf8HfbtY+0T3/uzY6A4uce4dhyWRZ89ZSl0CQasZ8NlH7qvZqVL0XkZpuJPW
yHlPdbi6m0ZRL3kLL3BtqPnRy2Dy1mrFXBkRKW4oel2h8flzaZYMNsMVxD/UeaD+FmDvAgydMJJD
4R7tbgG/X8fbgf+j1j6hwxZC80D33FwrUIkhuIln6T9DZ6ma2O/npJA8sY66LkEyoEpLRj0LK18r
rKKxAtSWCox4wguObYySsRHdJHYI4ETnqfTT/6PSfzd5V+neUui73NIqGBZD/Cz8QtuvwhAETfhZ
mv2qkKoeTK6tOPB/VMIIEQiuT98xA5Rey36ecKaXsg3tJc6jRzyTK96SNOyn4Sa6fDlwMkmnewW4
XYfH2DhMdhboEzh5Q66LkEaxSYiGemFDDQA26LN9NOEswSQ5mFj8pvMlbpcacOSFHKeYke01OTGu
l0qwzBuCmoECBPXQ1V3xyeN0xJJpVbkDmilZqOe22S8bcI8TQkiBtBn7PF/w9EuKoQH4bFwHc7wa
9AS98vRMSMs4Qp8H0rA2SEUMYxcZMBFoiO9SSPPMnv/cW1lZaeHeA0SCIE+beO5FoI3HLW6WnqPI
jZdakAiueFMJJcVzxgxuRchHlqm6vmFqBfZ/fne1s+gShaX/iXJpD7xCHKbzpRiiNxnoQgz3Q9QR
y6RQcnCp7ivvYWMLusL+qHjc39S3GApmJdc1YzOr38imrL2uNRNQBgyMpEdjX6dBHSdKwoXL4Mlm
UsCS79UpBvlOA+7dJUlXmiUZVoVeGjPfpnG8mo+BVxOexK9ikb/QX1uOLCk5ayaL2npmqD27BBOe
/AHldbQTUY+/sjRMPIDbFqN8q/nFPmjujet5mBbLyOtuZs5elgVUMSA4Gydowua4aW10oLf+Tnpr
5xpWXHuBMAejV5ZDuWSCBAU5MepVdyJOnVEfA0/ci4O4iLLDO1fsgGMcHvx9FXzGZFwcBNh/A8P1
3s6wx+PmG6Y/TbUQodSgy9sSEiw2QnRWzYsKZPkEH2kVvnGy7eEQMOaGY7V3GOnUToPuhL/POWwH
HQllrN1FnUFOtFFb4/MYe/BDRPaelq5p15E+trgzg02/QDssw0d54V/F+Wdz/75ZXdzBr0novuVg
w9RGjV/EV9oDYcjf6DlhcbURriQ1mxehcUacfH97Hd+6h72h5b1QJ17Kvyvo0FcFsWeiakwGWWY6
V16KwQ7g58yjlf0jKOKAE/8m9BlW0Rz052CKOTJ3IxWMyQ8EfzEXzFshWa1Af3nLRoSqxr/HIuOP
+RXleNO8dCHlbbvIZ4oU0yBBMWX86GDUDtg5k9n8Dl0GWKRjojaw3vYYmIKx/CjpDmVknw1vQs9a
idfih195js+sdi2IG6q1EBw60uGTndZAJpgyX3DhYIB/NNO1edF2MQxyXvVXC/42nRd3sAH4a9c0
9IDkCh7Siq3wu80MO+pt27fFrFnxdZ9fGmTCigBRiCvVx+xLEVlhGJiaxI2O6kdimmgGakaQg1ML
53jkCecdM8sGvZhHd/ybznewSD5V9JzMnKy/1LJ4RHGng633Db7lvCeI4mWfh60FX3kFi0ckckpL
jOSErSzIJK70XsyoG80ZSaBuJP0y+rCWDuJ0hS8tpL95HmpA5gibkZsE8uxz5M+T0epCNk06zdF/
fhnkbbSqrfRjbOT3xdNXGygIPsdcBw3olJcHSEyY0cM4v3Revz+LoIF6jNZpnYLPBU4geHyjc4j3
WHEgtUzgTkIcldHmz0nMut3+V9GerEaxJAgcqe9DbxyIzcnCeDvLm+oSynnKtjIlrEKiXyqfK1VC
rrb8BMB27IP7DgIfi9Czfy4p0T3nw/EeOB63zz5A2xt4eAn9V4iiG1Qa8oad2iJvlznNFZ7ywBy8
2cKO0ajMIKnNJuAP19y0nKgzkf+Df2LPZRhVAHx1BIVZMbOe/jodXHqpD5Fri16OcLLTLK9kvrPm
HhO/t35UiNzvFZE/2xZFKLXeeb62zgM1TaxTHRtyPEoGmjhu82wciqFFMag454PLjf+GYufc043Y
CSlB5AmaUqHcxEySVUDU/BfMgaEcqZc6rsZMFFT5jzvEHcnIXKpar4fNzuR/GPxZe8KWcyWjOSbQ
ZAxp9LQbxU+FYnJtUM1NpsJ+y2BAUfp7KkLuHQSyq5NJ92D680iUYwZFSNIiOMAK0SBrVskZwsyv
YXJAatQwBNsBS/93DPnd2aFGeoSecCQt2k/VVhG5Y0wWJlHuK4Uf1Cq1dnTa2EAN4I7LgbEFY8ks
FI6Etv8aTzYv3wD6F6yGnLjTxBat7w4m4cA5gby3zxzJzNLa99F04bqMlSjUa7iFdxGvIYGnOAV8
aUH0/s97DDXYVrDBuM97awQlUoPQYMTPjkHGCWSUK3OuU6ly3W6bLnyEEHbXbzv7RPJLZ1Zg9EN4
EyXrI0Cjah6hjLHyWyKlqq9dNe8FOxqFb/2Ki+kPLDKhWmSEKa5YhQ971xQGe0nbXIm/Srl1Pb+Q
b+LEIUUkPw9P/1pOgGR1W5fJgWJqLxDYJ9IKAqIkys27iVCM90804b6HeT+zJcqUF7OSuGDazPDF
iZ+cpXbDG76qOPnMNm5mzTiNJ2P7WS5wCSATRpj7vPMo+90vAMODguHCsiK9i1j61QVStNJqCSOp
g247lzTQKp9ffW6DtXcXVLqgsdZhOyBfLC7BjT8rOmQrM2Wd5C+K8fl2Pr5gYekI/1usAVLzRBP0
yLezeYxhcuFgJL1SO6kdPSFlx8EjRZRsQwOGvr+iH8GRbkrhk1FD5pB8QN37Y8NFbLRIVB1sANaN
xcQGeZptR7DguOY8KO9mlEIm8YlzewfiTgMbizaWQgmUctu8K2pAG6MnGzwaAJtYdQNaozqgieJc
gtn05f9UcaG/fm83Ghq3RNp+plb6GqiN0Aq7KsoYVkgQV8PhFl4fUFEncG1nTwKcMnm26BpNj/ad
hkHcG1g6WjhrZtgz0r3y3Kqu5DeAqYW9DkNV35s8C3yuYvjFpfRLAmuw+auXiNwhWlFfKwvE+ACu
crQia/ajo3b7/fUT0grH1jlmcHucfbYNbsFKUFmdtqjlqp55L3Cm0LekP8QF4Fi1bR079kjGZKmJ
Yl0y4itusPW3h4tGFhOodOwBJGrRfk/8LiATY1yVkJ3jf/sJOXfqMqoO79dc2mu0oGUzt0YewaH+
ixF3GssNaaUbwIKLIg87e8+Pm2Cnrxx8OmFTNOokcQt5NnWrkMimZle4fR2tADua0OerfkWLcEdm
oyisDu6i9s+dyWrFNFZKRONsXGfRJKpvPRSuI2sSQiQiX469PI+WjjAhf5/yb/Wpkn+MSPLTY6Pz
ys0+CTGBLQyizMCM3Krl2eMkbjAKIJkEAFc5eXLDq0hakZUdI4tfcFC4NPsBIXZl2Z7fqX74f+T3
TcsFD/CZY/Z3GJWHw72bky0pUdma26EAZj+JCtwH1M4c+BSkVemrdGWIW4Xut9PSJJl+7X4MezvW
HeVQlhMS/XoRhdg4Q2OVoMdhmHVD25UxEav5oahR72PdQREaiVqjfZ9b7w0qAwBQFbdrCbC5ozcU
iWzE1kKdtM0xCmIug/tTQwpuRAUExfZA5xTXTRASGcCrPpkyzTocVCHcEu7pxhGghfL/zaomeXLJ
5lm33Dzy/HBSlYhVd5RRkcQNera81Xi600v6yeoVfYFRmFZBPD54PdbZiIwvOxLX1SW99atxlKcH
SXTmCPv96C0S3gP1UNAibpwd/weJbtOSQRrFUFovdnyw25etLoaKDJaFuKpeY0OHRyiBv9z7+uZG
LKxeDm9c9rJYvLjpV6eIERG6EgBys2oViYI0+QROy0BO2hnYwGXONrbJWAbCjOqcNuDWFGXXqCKD
o+50smGlo7+mQVw6n8MdqaAgNrKdShJB9Jq9prBgnEgw87LWLXN9wNSn3sllpg8bGm1R2acBITtA
lT80UmNJUq4EY5D2j2ht4HqppFCf2qbpX7TQ4MenZELeYHSmGdcbkgICHT8aC7+d6PILZLtwxQ9Q
Nh59gU4u+QoMyLPeZFl5UqZYctV+Wy6XcA633JBUW+aIN6uhSrhmw96ehcJQLQoaHEL7mXLlDESs
8wlqg/P/1HsMq6fXRCAAhtir9DzyS8YXUAwX1edv8cm56UnGbPcClomuQd6VOllhg3PZ0s7VE4hd
pcJzU1hbHCddtGRzdRi/M2VE7c7nOi2JinLHsRiIoRdoG4yfbHnZVuTp8KOLY5hMkiNyv2Ikp5MI
NynKjQ/NdazJdYs3/V0p/TDmSq+nYezFgzirhIlR8WQ+PESEI2U0GYqwKPpTwKLM8yZkRUFCSIGU
PxejkZI/jEx4eq8VBgKijIT4UL7OL9REzSnb2iJP6t3VyjtwEb2FJqNQyRuhoTYZoARgrrfsfpdL
ZjE2pUnSAoEdjbHH0CllgVaQrKyDHYY7C8mvm4ENg76Vfw79ftb7IROmMok0U/QXA6JhxD8Ii7+p
u5ivjc4fBd/JXV0zPDlXS7BJxVmTljpSt/LUgiRU4gcqRzGwPhgL3UL+qRTJua4DDbc9vpWwY93i
bkb0B8ad9VtlD8TiQJVTFwrmxV/qem7kZ5PE3SBCN3cKfen+w8iB8nqgF456i21NH+zELTWdSzj8
GKX8IvUXRn3qHbdslUsQzgP5PPQXBhG6XQoVBWwQpPIMyGCZLyE1rx3KXW8zyxjww44cxH6F9lDV
LuXYGlkOgG3OiLN48mkJgh836L85VE1gV1MsHs/kkuQqzEj0jHlJROVAh54/F6Ot13eRCnE6SRkI
Fzcj+e6TW4J46OgJuR+Vs3mrYGE+YtbeTBdUFpcX+lhR9GOZApqI3rDm1zyMREdhqEEz9p80VW23
D9hxWlCBf6I9RgPmQbAysuEax8xSY/5Iq6JaXPm59EIyK1XSpF5c9/bgCQUnXzdfAFWXq4ixGnwJ
sL/c8tS52zpIZcBe9VippS0Y9eEZJ2duaxJpNjx/4PyeJGJD6PNM3Jg08a9TPzMmmW+d+UY6GlqD
gogrFrW4A2nI00Zx2pbjwnlzbIggnkBo7EtcfidjcQXjiEMkuMJwNL67t+qMmtQBt3SC40HXV77Z
vTqrWEuoldRpdAxqjVJTEhSMPZ8+Yy3QERnYwtqBEjdtkhJInmKKDdJTrxoPOab0yRZYPenT2xws
Ki46PomK9YCnFMLPOp/kcwFcoJnlmTpNZuBOCIEJE6+e4kDWSsvbFh+UAgaNugGkA/Bn7I/PHXli
zE5KEeqd5ZvF2m4bNgcbVi6Lcb5TRVU0qu2F0Cg0PupqIhXVdUtKDxFAp598dU0uPj7klHp7axna
JxdROhsNJcdEIhp7CWq6KAXkjt/SrDd9osPWI10RzNYpgojX61yqUo+R2/n6Lsa4QzvoS7SABN8t
TGsp3ZZP6VfCrBdQGvzA594xRbc1Y6VqL3BplSVt++OZL4c28ioNWCFK93Q/UetCQnqQCbL040Am
sYh4mNe67+yBTrDw9v+pjSwvsv4f14jBsi+LNsoxVIBQco6PAganw3YqZf0Urxdn/pLscZxg0ode
YofdgaFH+vVv3N23UP+sB08+vbOoSukWJfwKQrK3cKQoPFAftXPGdapnQ/Ul2ePljNLw/wDdAkVS
bsCXScMVBIgxFPX6u52mkqYKFbGJ/ZqeoFIKAGEyBsHL5AyvYglbW32xbeBkmkjE0bx49k1TlhTf
57tEWXxzVuN/1QqpYL13mL6SUz8le5+gcxPzDLNW11uWJG2DAkfTqEUWunf63pi1R4SAYsRIjYkm
don4jEFI0AoRP9+CGISH5ieaO0s0Ea0ScYbvsYUndcGwiNHURGtbGgjV8loPpJzMUHea/4WXgM6a
ajefF5LQqMf5XT+h5sAwSsqHmXDUHoU35Z5BTsKXdiy0LfYwE4spy/zl6HxAqDF4z7Plb2uvDBj3
s02Oy1IiVpt1tswztKLBDIx8j8GhSWLglNvmZhMI4hJzwrxdi1b8xDzr3thgzf6fDOKgkZa1+7CK
t810F7NgZLrQcnoEbeh0ba+dFLwCPmon4VLMre6BqP2s9mUWbpMabeexgVliCTmpGeBeJfCxxHXX
9/eIwFuJue3dVnP7k+Mv/POcw0ypNTLNzgGhyqBfgMnTz3Mn37Wbu6fQEGU1654AogKsMPw7iDw/
TSoz5HyA4HcgQFx/sgYGZRPVByzPPqn/jZa9gObI/1JEnTd9SshphP6DAbZ5s6VcP1BWUGM7COBK
wF5hwEB5uoe9Skk6b0YajU8vfCj9dyTCXLkScwoRAO4rzsmEGpSeR83hKMuGurMOy7QMvw4h2gbZ
Fi1xwnhuLqpf3hOrbeZkljAtaWxSqEDPF/O+F/3+0bJNR2KeSiITxJxI6Ep7BA4ZVJCtnni+/HKb
90tzTznAVI1ToMpjpLl/u2ArfSBUnkyJ7OTidwC8EP2MoGtl/1RupBObflr3gh3GWqR2i60aIh0f
fozNbtiiS2TX79RLS3plr+BQDKaW2FBVjdzff1VwyVFbp7gVI3h3+P1hs2dXpJs4AQBVrkZMWKS/
CyyHFl49EltUtaz6TgeVmJNEpKAu+K1EgRY6Mr17u2X7X6cvcZabmluhGk6pP0smYEntVNqqwPK0
58a5X1aHVv8fTAqP7TznQxhLw087oR1a3FyOiP9hfPjb+zmA6zHfEQlqxOZN9bpHV+AYrqJ98/i7
vxtuamxZQdch7QQsbQCuTVpdSxLtp8F9idKvSVmPvnSoMCn4E8UWWm/0sI5KYqNXXh60eVbrc1pX
9bVEzJ7vs9gK7Lm0jPfI3pD5/gOtM4yO4QbseCrcBFE6YOdQKarPRTQf4tWaKggHrBwSQD1reQQi
Qw0CK7pJEi7yB9tu224yg+x20w5ozOBrFs8G47VlyOFsmmzY2bhuTXbvvsduMjQiQv0NoQ1PQYOK
AUycbtcsnZb4Qw1t0ZEygjxzX4YOeR5sZbhnb68GkbIzJuqWK/rPert0512b5rTFk2S9ur5c2SDU
SDDz6DlUkGLi55rWZhZeSk1pyxS7wMpYl8xeTKN4nZA10i9kGtRL0VQq0jy3DDaq5d16nBpQQHI/
lwdtT1hCB8lABRr6xGXf3a2I8An2tUiOOqhF+O9wBnpLP+HFe/V3poN9VoRSOfyK2V8++NTl+3g3
Q3+Zi3GLcbew1Inedfy3DW013RjrmkYOblZeSI7ARAXvaEpeuWBqGHkGzk78MkA/Hvoe0ETeQ3ZA
26m30B38CPe8K1/iPWJzvGchH9tq3vV/u57tyOMrhJP+C8KpqRGON8E3VOOGFZti3A+DhKmY3igV
qOj0bsY+TsVeCxX66O0vnJhTF1TDPg3WIAEVjIprM0kOeKnjMbIoOijWSBlGFBNurSqgiaZX/o29
LelWMezakdcsCx7i5VnnQ+1oYT8TNHoxvU2jzBTvvbDjYgCPkqGCzH0vDKupBxI6Xzhy++ZliNUi
PbiUnMpdMLTbMiQQjpNu46YBC0j/QmD1Ar+qpopZVl8kwxAZ4MUodnJDdWc5bqyyY8dA7XhQ1+Ga
5VOnGueILjqOv6OzuqpDYU3Wd/Ns3q9fay3IXxcIfCDZDJG1sXjssGI13rGngX13NcPwdY1pZ6KC
pJn6i9uFQD+8olrYeXvNilEIK1RezWdTKIjYI0wl0c9E25+s8g2uIsszTTejXb2UdbT4a11oUZMU
6Q46AwwjZH63YU3xyTuw8D26V/4ak6g5ITLs0feLVmRqrI8HCYrnIb0q08rLlcBNil8mJvQ7Q4nr
YH/w2STT9T5RE+kg2GU9f70vg0P90yLARHueAorLi79qfVFP1+12yOQ0Ad0NrbIVBY42sFy5EhHY
6H8+mxE8zTFXPTDY/6xcSma/1akdBjBW01+aWvzVF8/bzRc/7Fz9i3mxMhsH6ssFskLZVH0kH9YM
teXuLzU5jAiIu6ZS1lNjIuO8RDm7a0g18i8vcTe2xXsRXo9AUfPXrTqdTsAzd/zA0NEBpATb8H5O
Fr6kC++p6lSkVj6ajYzpjxV1Qhm0TrNV5oBkW3gt6bvF5l1S4bnkO+MB069J6BDQUKzBLlpI9G+u
US6O0bHSNKd77r8P3bRbCT6Db6c9C5KZSSjLE9Br9MU8aIulvhFb0XzmG7TaRHJUPuGFZnDrYJVx
+L0rQRgjgW8ylMKqbmK2rFlNAKreVDrphTq6MKi4JHwP2XRuAUS5M6X1MyTP5w3Nv1lwdgvzGXJR
SGNIIWQUeSyStDMNq1slCcGFBool4O/DYfvAMDWmOdNtvWuw5hWatx2+1Xx4QtqF/uEsNtGD4JWo
caWJ2MloGjDsn/aAmEJzcnWDrGVYkTDK3rYEDrn/Rz8Kg/KdtETKYUVYWIezdO5bcYCa49tmaWZQ
j8VI/kVvNf2wa5p8UHr+P8ydfybV+pM3gnmOL5OHOs7IcKfAuKmxdBVqYmCR9vB0Qe4ELx9vbWUL
I4Srt/DgKCTrK9M8ukhIE4JAYHooK+gEnR51WWU7frl/2ZyInmItZQls9pVQpaHoNvrXmh+NT1oG
eBu1TSOBfcAmcS1+gumSRHLmTe55ittUN+HfbMP1H8264PksArhhWO/sKBe+7s2pcMiJgoA/gyET
5FsZJttPqD0IuRk6bT6LX8lczu8k2c8Kz5/oaUBdNjjGqMSb7R6WLFbQjUgZTJGcvzMmmzGX7OtV
Fmb8wHa8mtmx7p7zkCnYe+03wC/ZibWWFTJStnPribQH/naw7rAZiMEUab9W9Jl1L+XtsoYVteJY
WDI0CfKj4LREYze4vNgVayJ+jtKK9ryC8wVsZK0uzqco3gV30EnSQaP9TgJRvtbV7wKmGviQyJpY
IZQCYEy/p+sv3WlEVS7ntULz9JjG4TT3bF5Da12/mxc35/xVvFYVdtgm0YNmuXN68B86Fi3dkXlO
FEQTUERVmEXpR+Myem1mNLQmyfM8Ml7a0KQ8hCo5xDLrlksFFjFsLQGLtO51om9td4vcHQcQpysu
NDzkx5PCmukhHE28X7u7qZCVlwEAzVGKOLPmZAIvIEUCTTOf3oIvxsGAy65OgKVb+zW/xq2fHZE6
AopcsMfrQMSzuJFOFEEcIBllwGnH2YFNsSftL8Re84xYm67gLfaMyHM+Nn+EgUfO8ukGvhSx03gr
WCe0Bv4doY1yRUyD9FPNmAisc1C11EMNJDC99gRzqABiCugCBvehJq0/6GqVGKqznVnSMPpweLFW
yKX2B6Y6C6W/05QYcBnBpsFAm+pcaGeubXLnXOZlXKrY514Ml7qmH86cI2pTmeWpf9m8XrS2BdHM
/02oCpLFuL4fhv0CvKTbFf4hncy58hkMJOcoibpi0lrGY58U2S6OXdTRYS3mVqlPhxfuzr6UGAKY
vZq6Xd51cK5NiVEUF7j2VCdnwfspYkOyE1hIGCKngyrjm/OIZ9T2rc3z2ymVnacAywobhl+s5bm0
fQIndh6gVmhHdT1+hM/IznclSiMeztiYDXWPQ6rDmwpKohOIFnAP6x2OAzrpLmUe1N3GQ2cOV28P
GIWS/OFcjDQEBxU5MYPtYYqH75YVFArVe7aKEjDjvzUum4dkMPl57GXAsxEBjC/3ucIjRKOeE0ur
2apJHPF43B3Acvljox5JoYDu56Tf2ulzksl8KQoB4zFyswKvdFzbZUTKS4yN/Ppa6J0FzOHfnB6g
wIndggla58ineJuc9xrrxyYKVEAEZ7C/nM5igCNYSn0i6mbU0ZY2KM3gaQ/upZ/tyQ57Kr2Jvf1F
O4RZssdV4dDthp4et2oaGLUtYyxBaNmi2lHR4rC7H7LgUMp8zevlbAM6HoRFMKp7MFsf9Yocbopq
8Uj14j/FKwz7s87DEdxHI0PYly1EY+aXRixqT8GKU/W592DbCVw3DJu4Kk8TMFCfvExlTHM+0Lzs
3lOwUN/b74gpo+PSzaVyu5AwA2GnRulQtTr00viYydm4Dz6V8wKo2wZUAUYmy3gbj/aiDCrnPezS
XgUJ1InohvC9ymukGno4uPxHrupsU78Hweueh/KP7ITsF9447As2rpF93RzYUtorHNwLLhwPPsCQ
35LPwLfxg0jk+HbshnA62puJ4Zmq4I5uPIyJ8jaPuZ7vf4VFgExo5RxnOCc+bUMWKNRk22KROqOY
xkv5CKSs7S7vW88ZP6dzdo8NL1DcZPhv7YoESlCA1gJi20Wf+IICFjsOtaz3DOMwBnxgW/L26JCn
a6jL3Tn/yMmg+kd7zyD/zRvU1EQdLK4QW+JPH7VKdbrM9fk6mu2lQa6EBNfImIgXvdVgqVJPza2f
/ISX/ygVefQnPYs/xe+QxwO8EvZX6GYYAtGUVwbFunEFvLPmFrxNl8zs9OSK+dld0p7Wg8LYYOwc
0FUfWojSZ11lIDWe2Tos0f+RBq16Oz8t07C+75owh6+TvV+YP0M7AQg3b90ab9N2rq175rNpgTe4
j+lJzr2ZLtMk3OAcc+4PC+KLb9N5nolYYZCy6D8e5k1COzoYjyUNGp90SZZr8xbN9H9U0StYdkne
3/n2W7+rvgfquVmRP0ZHXro7iQKVrhOGISodwpODZQoVkuTfdDAGDnrTStpB8eL6qzBqW04ACxfx
Wqakf2FzDQM2QUqb6LJZ8qeNBLO8IAm2gG0irvQxLdqvJAMn7PLwDje0c0gNm1upPaldxEVxqKI3
0W3a3hGgYbd/OoVjAKIeftKpBVpfjbc8IpcrP8HEfvAqvtSfmO2EGkEYpPX0DOQNu9iC9rGNV2we
0mg2im0werkwo5PIGNTeQVflvKepU9d0diaB+wsuWceZAQG4VjX5UH7R/N6KWWKayFXLY2frm5Ig
V4AjKg4q//Edo5cjDZg1mRH+GwEAhuP3ogPcuqAnCbWFfKNznxlX41TOlA3Q2k0ZbLLwZ8llIP/e
Tz612tuLms5w7TPn4vigyh/Zo2qr7MNCxEwBgN4zvI9C+UTBU2jgYicDp4g8qEirAVYnvulB28NM
n2ihWqWQS70dTqZiGPLnsqlS3i/S3LoQfjRICoGG59NhXy/Y5wokx3I3vNAd34jf6Cj5uDchNJZl
KB0WYiz7GTZtIHdu4l28DUbjMF+K5Y9Ebg0bIMDBDDI0G3pzy57kRWH9f0Kt5QVMIB+2TdR4lvj+
Hy+2ArlTV+kUctJj1Jnd20W4z73I4PVwLixAAWa3fhpQ3YijLcDnyqo1RPlpBaJI278nZRfJT7ic
YFwNgFbjDbxnUwJNXGxc6DfSZgLvxDmc7Ar49DptFtiQggBKxHePwL/je+hOiNQrVLZqWFFuE2zO
2DQWYRN19hsj6ZWvemp5imb3Wjr5BFAK2AJV0+4pXpHanIeaBig/23d56SC7tOvTl+twyX/uqnmj
M00WDF8R7VuUVemVZ7w1Og67AH4vD/ISnn1LCQwCW+IAE5sbqXAQVGcUzqAuMsq04cnXZztXjM4S
XqwOYOqvilKrtvekelPX4AyiWZeLo5S0LDpbncaH9JnSvs1lPIiK8l8bBHp0MywI3Styud+cWXWt
WAz1vUMqxwgohWgRyFA5XRZDAU9U//at0AN+5Xyh2Ny9ADEzWB8AgKSn5iqoNdMvlBt23xa87Et/
riTSoChSof/CDrTFAxr6W7hcpnzYIOwK4KugS37B3vh1EdG1BfhT7YjXi8qKTAccww7AkBE8MNHD
Nt93FgJAtbCUSbjqmopyT5E6EbJlAr74TmjUJCIBVNGv6mqYR6utHOnBQ8pal3yXkTzllr5WhWnh
X7bzmpbniIXe6C46YGgpySTdTQqq1yJOzYTUKVW9SMyXVgP8t6L+3O22pG0JXngQfcvMD5kDPjpd
UYD5enEWmiek2fbgXjGXwhxHlJIAnei/KXdFRcaBBNZJ99UBLiuM18WjHv5h4qr1h3NdaASPKoyw
K+l3N7XZrB4OIjwAH4t6lTxrJpNx1C74+3wsF/n0MYB1F6P6bWyHVe75mcVGANCimh+pX12hWIDF
IoaG9U3tiQbS4nhqg+805bIrXCPARrS5roTcrT82V8e2W7k/shpl4CoJECuvcrQoHX4OJDYLHU5r
9CO7wHovhWcf+iMzgpHNgy5r6h9hPTAHsmQBilhNPM0lUYwUF4xhELOdpPJMBw5ST07UN1ko1vai
pRqNeZ1R+oERClVzsciFXWWjK03xPAn8Vl0SnlA12tUCz3ZQ1lnMJ+sjb66iirn2amnKhE76SnLz
fRc6prAsLxe+7hPvUVZ5MnCA9PLSwfnLv/XbZleYJhwECaH6qqP6BdDyvMFa/hmyN0RWU/7PB0Ob
XDrUGfErHZrl2MFa58zyc3red4O8JKAPVRoeCfti8XT09/VzSnPbRsPT6WY0/9RmGXPoaFT6TqwX
PIxT8g8Oiawhssqe9+8jUGVQaHMbk529fJMNBxvGiUsKJvHmPPHWYs2TKBG3sEqUaFXOpBt0uefw
CHg+aMf/5exguqLFQCXiKecpPlXefM/WjBa9bhn5xo4W7K7hw/u6IedAbGFu3oJo5GjVY87ySlsA
r5XAG6xzwFtxUic7pqbuo8NDMbeN/TRTNt3dwpSbjzfdw5bysajjuLY8QR3zqhOTC6zGDya9hLGt
8kHQR4iVcfBxzGZCffI/6Xk+gfgYxXWbPPD1XQVcly03/GYVUQaS+GrWbyL+vTCoit2HVmnvb/Jj
lACk9IacoOiWmQwBgkh8vqsD1EBy+3JeeUW34Lh7iOtgPUyHdwAYQdtfeopmAM+KAbGBS1dzr9xe
3SsKAXm4z738CO9tmZScESPZXh3l5rhbq5b81quiZ1I36KAuh/3zlkW5BQeIO7yeZcU6+qx18t8/
HNuZqojxGBfkiy561p+XLHQcU5dlbjggxGCsxxyZSo59SB6KgiXaUT7XJHLL07Zoa695oIrSd6sk
DunZR3YFh/Zqa4hF0L2srsLBCMf0R8AwsQ/fQQ8HBgr27tH4heHM4dzL9WgBzA2MYfy2rnTKEamo
LfZMP1rddiFuMWPKeAF0v2AADIAra0FmiOn1iPwz2cFJebuJn5467Slb4gZvYfP+TUCvyfmJNgh7
dXe63esjLdXM1o5jsWz3bDu9j37VYLN6L//s6lfhuhomyyAJqM7XZlQA2IR03rgkZYMGApngJ+Gk
RVUgGLKsp9h4fXl5ccsn5BJWDcZSa5tO6EavY2HgDtEGARu5S+m/CckytPzzpTksRPR3uy704MQp
gQOHdVPbVmFoYkhb09FNE3s7k5aAj2jFfSI2+Ywh6MmFEhg231w/3Cujah60LJT/6c45NcyyjMWg
QAPrS4LNgRksNKguP8Jc80Y/u1Kn2Temvs4ACyi6HfkIWbzBx04HIOfOaWz92Rpsa/NnA69gLiBb
jojiPfPOU+9Hl7h0aIg/meRwnQ6FZppK65Lsq3K4/bNfETRygVI82EnJ78EAKs21lfkYzAZO8OPr
YfpFfL0EBqp/bqxs2Egmw2S4EA+/qRrwlamXD4csCVtfeQFLnKU45rtHgJE3SnSY5r6pC2C+9QxC
khe4KDhIGjU4b8/wJX47u5EJB7zI+ZHzxtzc/9z36ufB6IsFttb93AQXbodQyl6rJZOQVi+KcOsM
/oHjE5B0giepKIHGyKhqpD0TqeLd4+X2zfazQ+1xadCXo4fbsPyQqpXgDJBSko/LNRa2+zN0gkkz
uPJdWL8Bj0rirWmjGJvuhkR1/rh7Fe8rS3Fjt87lBYv+Xfm1yJuNy4/cfUQS6g/KGWIS2Nn7XpdA
nn+e1WndW67AxVhZYmuNsx1cVaXd8vnKbvtVUcK7tTEDhigasmlUMOqb8JGUUrXQlfe5RCncShY8
/cCPyeOmd79KXo/tOAF0tzdEQWfK3KI71zNY0lCvQFDiUmYBqSuX7CFxLWs6gRbhGHqWaxBK7dvN
P/k3SArIXI1htfwFmOfrUVtKhrBcoKl21E9u5Ej0QLrQnB6W+WCgkev9WLnIEShXjG6aOLrvbnIu
zZ2dk1aaLUHIKeC6xtjUmXX8JJ9Xp/sMnhlKXhsiquwpUvp8kREOmyZin3LsU5lS4JfFZ9EiV4Sq
VZgOjAav4XoHQ1KOr+j62RahbTMEvh30PEgRXEkoNaD73NPpvlxqHDZ6oU3MWArxUpeXG5US9SVc
9K8p/INLYTLJuYrvFMpAimHJ0vGJO7n96UnI+dNJH1haK3+KlG/SBwtNS1iK3E4YWFezDNADte+a
bywmIEJ13GIWGoC6jh/CNMFDmBRMsWi2oMt1Oz/4r+mVUKOnRGGR+2UqFiMd8wssRVV51zm2/kGN
3RZDIpfo2NrJ5TqJLz8KENdSTHt5V/ky1+PMYlRpquQ/Y9aJ/58lqM7OATDSuRKIiBapQ7ngfBOq
mZt41m5CExmHDGWIH4Y43lW+d5W5mSj9Q58mR8rJEdH2NaWkjQsXWyMxkzUYipwmo4o4Xq+kqcxt
7pL0tBY5IFAbFh5dFNLUaXGzhBjDUSjqXz/kvpnIMsJdHi7s+uI/WcFApkG93O4QlQfqStIpzq/O
EPFzkOroLYwQl9WVjmjav+eLBug2h+Y5F0zYCaUcSSCg1PQuSl9qbbeFGcyAQ0/LTLacEDONX3sX
vWV+yFAybsBrMAIEY0Xm8CrW6u6tKU2xJtmpcJCKYViK5uCtIDeydF4crHYdLQX6U16U5f6B7iom
xsruKgc6NMJnW+F8iiwJB2QcDEgqBi95QaRFP7LpuT+1vThjeS3qODuCxrRmjVc06HJmj8zWhULH
Nsv3r66AWI6GpyJcVdpi2uS9UUDa8k0IctFs45ou06lp9z5+OHqjEAannBbgLdWddLLuO3XwzhVj
tVR+hYvFXieTuW7JXMCEow49/98PoRzWPW8WWhOChHV/IPv4jEdulW1NEpCSqHYhk4tXj7RF6Nz4
0pXomoTOkGsWYldW4jJXUoeccH6CbDMjRwfTbN+RYiKCqsieuh0OMaOM2zZqyWsBUKF8uJ4B3i8T
DCuFK7BMs/6LdnsYfnUT6a4EY6xXhBBTZZJvHRI9+FwyZvXo9cEg04hhpOp2LdFAUsmWM/4xPoBN
PIi+TemaC9lPfB1mncgmeXZpxih7GWi7OG9JEqBcc1WdKGBM/fZG4EdMWFycipRgg24U8HexZblq
A1gBzE6WMpCzkt6pK8E6CYmBGTyDxKeNSCIchXNacfYMmRLKsp9qygvbA8gvOJ2EkyuPiN+cW8Yq
QnGqd8VAWtcDKA5YegJ8THNLoQTdqlQxGcBOo+u69ODdlDKL/i2xwkAg5C/UJou+v3sg5ffaZblb
/1nKwo9ItjnLCT3jVgGGVXp0rfOZMuTrv+7xgj0MCJpuXtM1kxJcLki/WJZRFrtNKuT1hmYCOFh5
tmpUvAPsslhFdJsda9r3cdhjfYkkrJ4lUAtEj3uGzqGVOgQ9z5K3xJwbvJ3ooKiV7cZaIxC/iwd6
yUudBHuqUeClMLJApj7JsrP//BM69cbj33NDyGlEDOZzeHUOpp3BuZqEG3+P5tNvq6F1MNQZUlOM
64k4yS8yFXJ78MbSgIwgYPIcROtdss2QfEW/OhaBl+mJJu+LKTWqcEW78+j0sPFBEkN5kjj8lSXK
Z+YCDQ0CEZU6EKHW/aDK/81XBLgKkv+h684esTukU0WKm/+z4LrP8UarhJcwWB8UIGHlQt54zs9M
QWUfffeOGvbkTkK6EVcVT3hOI7zlUQ8+wAzmzqmhjne3CMA4TOnPYPK4LzRe35X+ob4c9oIJN/or
GqICHzRAbT//umlDkwePr7mHs609JSuRZMTVedY1JLmIYuIWlclM7PMnDrqlZqHi0LmTdd6zpM08
DCL6u6nX8VWcfzXjLHEqAkt5lLkwYSoRbTLdsZYGtLyYyQiOLoLiQPi8X1BhPaRFqvY2wktL2Uwm
91GlBTDVTqGVZWXbexrtBhxfclPzEUH451CyKeoyWPyUAjPj0TrsP2VX0Lbq7aCXECDXes9J6Mta
iuoekUHvA2ez6IQ3DMHSdENuJYM5wjfcF3GQFobNtZO5GfKqPQGJB/tZWbJnd14UKo7ZRWYteCds
uzJ+snK2VTMnGyWRgWl0qYZJYxd3kvhOD6KtajYiXqtVrrqMT3ywmNZ9CZjZArA/NEoINnbWHL8m
dQ1iroEeTIz9gThxrEaNs3cf6YBcHiJq2DIQ/eBDT0KkdhD9wOKWDnwvwccwO0t20rjYSPs4bWSp
BErsnH68nMp1EPEP/LKw4UxxoK1ETRVLM7uFGQeZQFB3LBA1th3RBG7GtVQmMuxSKVHPA+59wW/K
o/KdNYOga5hCkHCXtvCaBoKNFaIzbPm5ppNTFz1+QRkjRSUZKj2la2Tine6OlgEXy7a5NMwZC9G8
SDDs+YADFY55DRmNjqYLFpBA77atqawXIP8LDlp3eccoz5LmyruZ6j1fFb9CjSt75Cun4PHiCByv
LmomCd9Zy7CVV8th3DO0UYUSK0ZuoH1dcATzTDnB+nCuwyyOxBaUdGKTqKXDe6WY2eRd/6gSjjtj
DHpNn5pw5xPGkYcWmfZ6fhhpw6JicenG1RzBvFrMuqy2u5lzKOrERRhYSUW+PJ2gMN607YVYOE65
22RnjgqjBE/du7u/nHMMW8BtQGUKKlvv1wbeN97q0NFAc0sSm0wq9QL3yzHQhrPlCPDaB2FSadLS
30RhSgZhPGv572GCgFtw5M2Lk3E/31PcglN1wzOmiExnZ/Q/MLRxEUdcKzsuEM3YZ0eeZ6jlWjKW
nUjwORQZI7M20WtdGYmL7QmQ0XIevwWr5X683h3dcQwpStwZrswHkBRymAmzO0UKzyCy25Qf7af9
1MYNxcY32LciXoTHyyf+PFG8M9bj3JRTPY96vD3SmHVZszjw21E1Q+nZuZ/LfqVwJFLSsuxlStSA
p3lhSmosbzfIK4AfsauKmNV2jPnasLEpETdNv/uIlOoEcruJE90TbSmQAMGeO58EPWnRBlpxLT2L
ImQWX9C63BLo6uoBptespk6F4UyK+XwpYfiZFb4vsmgi16X11O/g87RhWmtMEeZtkOCeyJIADWyA
FYAhFdEXkCNdP0idGrzCjfKIrbf9zPYM3bEIvwx/tfoF38r+OpFg5OXNrzIcX2ozJTJBjY5t/yvu
j10I2gxaKJArPyhbe+p/V3QsH9R0RZXD5Pq68jyMVfEEje4d59Fc3BLws7Dwdrl3O2d2xAt+6LAB
plq1BDZmg1NTIHg62hVSC1+hN4kcNeaXj3KfJLcshbGhZAh91rGE2S+mgmc4l/Itv4/kvo7M4eXW
3b1A1umRQnRzWZU3QMOJTFpeonUzsd/XVCDOTFz09+adMpI9WPegTYsAkl9R9cbZgXgvHGhQYt2o
eIAhKgZUxs4f7G0Y2tjk9FaXq1xiANfwfRv7j3P3iRtjkvwnpv+lZ/T5/jlFr55d5kSDuQpX8wfE
P3NGge4u8uj6QBr6eXn5YJXYVX38WRcyxUrUMAylPD/ubx0UVQlYi3vIZrjvsyqSaYU1zVaey47S
9IqmzBmPbd99LdXMC1NUG9Uhpb+ujigyILTd8ez2JI34U41O5+FCtkAKSXwOJ7U4sPiX4TyE1Gqf
WetNdx5JJ1+vbUAeiXUIRu2AGJ5KFNUWZsVDBCOy/H22igelxW5y/Avlv3UrI/+RptNpI60Ko6Tc
+NAcGhzFQ7+8C/iHCTA7JGX9ZKarEyJxaZZdB+SzBVzoLYwMGSO6jE4FPw+iTq29yS9o8JzbllH8
TfNLCm/cbEEhmMIABvvF/UkbDApvhQdjEVj6qdv6qpnjZNNXtikZh7L9LudZcuJJqXmxQj0IRMg8
5Rlfob5lBiKwP525m1pXrEuvl3QeDUvTmoBELv+fv8hIHOqQtjRbbsnVjmSCfzZc+E//LL1d2BcO
vOK4wjBoYeAtdN6MTVEem9dOj3YxhpGl2KOtLBflBOpOcNv7Hh7sFjpIuJZKPWM7vUAihJPWrxXD
lxKzCInrqc2He+yxKL2nU2gXWN5Truhcvq+Jqh+a39e40tVFfzTLF8D0pzXePilI/f/fEdpKebmG
hE5biYG9FHpkFXIEyVzDpwWE9ZeC1HwtSIwSoeMve4Es3fFCCEZtFZRHZ0dLygLsZjRVEwA7Gd62
wb1bMQeOHytdwyVmB0m1bYuwisRQJBnM4em6i/yZzU/9XYEuw0kdD+OU2tIFLlyi7t1OW0UW4zE8
HlnTFzXXym2abx0IbpDv5Pn4aYzc+kq+N6i181KbTAEtvaOjzPEyHXev++MiFa8d+OlMU+Ytr0R5
aLo92QBn7zg3XLaIkwZLi0cbhyCjPWgzuXb9uTf9RM52viDYVZhvW8qJ/oTOyNBdYZlcL/X8iIYu
ogQVSGu62tWAQMkYjQLahiLFqodnfAld4DzU+0izn2FOnkK6DjHZYcL2FwyI/n6WMdhCSPukBBCG
IcyQfONb76lbfaD/Hq5vh67EkFT0zXD9pGarNWBDLE64rRp8/Ctk2n/vgdcVghzuqLJcSNJ35brE
62v97CGFC24LbkPoaSC8jAAlCqUz9/OnHpshpAwWfzAUoejADnrm9GtxyDcofOIQwyoffScyeAuf
qFrhB49OmZbyzOMsDd6LWOMwaYLPyfE8wI75JrBeJj2JFLnVp78nEgZrQHRHOOBPaG5ZWWQlC4dt
mLNjvH1uiQXdBxKDowVeBmmRmfJq//v3lqM9O9kYaTRe8s9CNn3M0ckdH/8k+vckw1HZ8+dYYEz+
Xqdar8A2R3a1Kf9/GZgfXB6vNuD6PQcJyz4BZ30zFhwq9iCW91fDt52HjorSq24Z0V5msk/DeZXE
wesghMeo4WbUr5pVTf3reSKBvil/RtF5n/d2Pirp8vSTy7rzydv889U746tgU1b4MGlLUfa6e9BQ
HVXDNi3j93h9OQ+++KZznASrXxSUVyvluWScSfjhokTE88f8QSkfIkoN9oYnwgsAODTXnlI2Iny2
VWxBwCEfCodq6G8BqbISvENM0yyl/lbw+RRqwzMvOzyFi8ogFHTmyl9R+maDE9KyxIBp+FJSGcQX
GAy0/Sj6dtrFi8Y+9ljOXrTi4iSnWGkqEETdVZGtU2j/Okuz50SIfeiJsR8esOeDR7w5i1b5fCqo
J9gD9DhMFV1bhaMBfzb8y4qfb91Cw9cKgfMM3z3KkBVf85uduWL5oUYEZyEarWXC+3VNmIitTL8O
EU89XXVRp7xAR+zAsW+17pjeGylK/QoIGjSY/ru0y+3keVfQPo0y4NjvnPjw7JlgR1Peab24SSMQ
uA1Gm1pq/lv3+IAavmADSpst30KkMe5skeAHd2iFe1qrKD2j0zPCy+GTu50tWllejeWTmFAsrIHO
XRz2Oz5k0xa061FeoKPMvXeINqbFkBoejYd407gi+HuQ+5kvONx3UHlxJ5JnheGPqMW14HF50zFq
5Hmv3GFRsbS64yOgQ9oIKiuJx2WqXrOKHW8AMKUgJwl9zQw9wlJ4ZesJp3/SCcslao2zpmIU6hfU
nb886+mWKrHlvpAZ1mR7tlSXvbh5dbn2cVpDRl/k+jJLV9MCN85mMLdOBOwW1ccjsGnCNvAVAP4O
IHzNp3Yu79qbSR+nI88RcbfdMODEXn4is8fje2BNZgZYplfHCK+p4SWZjDZeG6uW0dyRN/vJ6ehr
Qn45zY1xNtks8jVh6wS6DrFM56bD+LsaR14vkV/kM3Q8WesYjB4UoR0iIi53ISde6CBbihomkE+2
lATmqtqttOvmV1TcAVTFMZ5gTCC3/a7QhJDlhH7TzS9hrTNxd320DQPKtLnRz7Do3KVkUMqPapGI
Fcbgep1WyLmFZEYPGh1/Exv+MG1zYwF+6BVRktF3+Sk00fwdDmB+7DAvn0PSdVaL92nAK8wjzpEu
CkkshkzIS8wT0Qlku/SUS5e/xbggAgu6t6GYQyZOeQ6v2M16VYYp3v7UBpTkOwIhKeekfe3f9RfT
rerY9CHSy8MJh8sUXqxA+7lCcyZvOzUcNVQ40B+zewB0lQxU/uXKG9LuAUAG0VVM+4dhnP62ojEU
f6VgmXwkKqo8uGm1wDmkkkX/GsRhF9ONlPkXWvqJeDrpm7Hs+wLGbUt2MKE9DWTRjX5OzHKenirv
Lq90bLThUC+O7NXFCsn4JpXgXtDNJmm9gmN2Qu9EIM8frxCfkD5fzgGcLbafa7fdcD71G8BGNkNc
4OnQG3AfpnOMfXCOlkNYlh/bmfHy9kA5NKL7PP0ueoJy9dcpZZ1f8DQTTuv7evztyAD46hM6E1tl
eLe68ToGEOixJEY8s0d+vh587AS/zezpa/YCep3BH0ug+xsyjYPxZSy/RUuAOfdDzVAF9v5odHfF
u3k0XAlpQhi4pHVZqqz7ZHvS7mK0IHaDTvvkgaWC7H3EPaR+V36kqibP/QTbOcjH8YSzKSajUUi1
rpi3/umo2cnlz69dGK8ty9xhHkY0g1T+AouVaDjXWtZfG9AUJnm87C8lbLpWq5EjTiW2aAbgF5C/
q25Zhg19N4lEmTrPxHXrtXQWkkgiXUUVk6oJH/swjU8NkQMjXTccpGwqZG2ZPCUE0ti8HLO1j9/6
XIUI4RZMwAvoQ4SZ8aE+7v6JNm0rzPAXOJL7QfjUal5fpLjwW+fFTAU5hTw1jwXuiySIfmVqqCYa
vXZwIP1MkfIph3S13zbp7h3fg7CR/Evl9zwtNSL/DEann7NEmV8CQbEStgDprJIS+lsmKWbPK/xY
Sad5pTfx/UIw/OCzeUdbiCNkKOQtphGxqS4jNkOZOY5cplwu1brWzf8SvY0SLdZ8nLN3iT0v7FOu
tJZEdOmV3auZMNrwtA8/RQxPR6iF+s7MMfdCV2oDkki0dWN5omKPFxpnDGhKhSGimegs2Be0z4/7
DABiv8lxOk4DhdbuFl1GpGez+qr5Ve4MzAQvH2UZZT6S/qxLHiSlxTJLTjvI/JdDqxoL1cdhCFMC
zFfYnS1hPHGPrrc5F22sVsHTGcF+BEO0fRwFslBT8uVe97ip3BuRl9IGtily7vYarzBo+lmJHSvd
02SKd7B4ZNvSoGlRdrxkM3VcoZFTHpin37dn5VpC0sxC/TyIyb0vEMYNjgY33ldGMmy5jlfKKE4K
xqUCj6EPIPtb9OTtCsOI0klnMifaUCRMUBZE+lopKNQXHNCNyJWRTUYnM85nMC2AMHi7oYwafPTn
k/uOHABATZn9IKLiwcLwxWz5/WOyCe/NJLA1jNkXvnOO/sNRtwXnoiktXi9hYI1LoAue4+9q9Zgu
PFj8XzEcxE6ddUpBOKv6vQWR4cBRSaZ3OuGqr8BYVkDKPbOTXu5xlXySH7nxw+0+PuKgUUF4hUIZ
MxmSvRgImmWCqj3FkDMRPEOu101THnuIoes14RIN+hNBJyYo3psVXBhw5bCIw0DHzxXk9M6maQDj
VqLPuzjwuUfUHDjq+2U9bhDdVKtbMQTb6bakxE5wsByYKeSA5QIquwQspcNMQ9gdnkJz6OS8/6Td
mD01IC1MONaAdNa20C2ZZ6IzPQA+S4pnSVt9fnekrOUnv7waf7molEB2RBljPhbFgPnYkbjQbdq3
Z35PED6YiFjbnbM4BNwjXl3t44ZpgiLbsFTFcSJ6dzS3Lmry7TgOZPnDVb13tTmRs/MskKQQA1iD
EsLWSEZoKdJWRCLGk4rU8B1A2ZSFZOCmSvlcKIrLDtwEEaO9uLo02DvYtUqOYD6LhhCk32D28ZrI
b8BAxlQJCD6dtKy4vVn1OnsFQNQap2Z5rWaIivNE9HR1LSGJkaG8IM4LQtViby+MXok4NLal5PvH
Jm7e/gsE2POPayHrd9n3XBktjn/bZc/+3tN2MVpL22IRJJGmRz5mWOD+Kx85srARS3Z3Nk90XQrh
O/VpoQvnq3YyYLZfeDa9Spvphefk+sP6zxy++/a4jW9dciA/cYp+kCAnckSZYsq0xy86r93ZcOQq
KyuXmQixxmuU6W+jIof5dIXHHXQHQQ459eiu/Jz68gEkC1NUh1oCZiXKx/ajaVzWfgnKXwTTVQRL
ZQGLhbU6nhNfx8xW0B7+JXk9xqr+5hab/RiQlB66b5xa9DPoJSQ8o7pFppVT/CcTzL9OCokA8SwW
KOvsE3TwB2aU4OF8Fgh1S4gle1F6Zlv05SSK4C84rnv+VfvWpKR4X3HgJgYu+6aLapWS2bLSpJbY
0Qi+nb3xgYBunYGYGvJct7xxEILE747m8RCR89k3DRh/7W7L5LWwP93l8iaqW2wYP6fxJ3EPSC2E
i1qDtnFqyTy8sRQtBjE4vlCsbn+n+yWPNAG6COifORcMKhBJ6zZUghS7ZIJqEcNIyBSNzQyG4YBh
GLKIp2JSLz4+kVOyJMIoy9OeLIWQpqRZr4Wdl2zXTbIGKjb4K2nIG6rB+wHMxTg3Cf7zr955qW7y
NMwS08dp3q1ABz+9xazh5Q8Lyhyo+zN6pPYOsYrhGF7ckgt5+XfCgiOp8jXnN/X/ekVdokFLdoXj
QF2x3A8Xpndz2fCx6khaIsJv0cLluZAhtQP6RmmFtR0YxTKY/iAlCInZJNga4WRy32OvhmXQuBKR
OMqWWpd5RnsLi1oGsTMJGizvTlWHZ2psSJVn5KMdo4YyjhXZzVKdsCpmTTD1JGjsannfmLufxdOz
shPjXBiGX75XL/hsXNPJHEinyQp7wXAApneG9SiH9755QQ/p6jG6lU0mtB0x9cYVF9JTwIcQg6ZC
2Mg+mvKmLXZED3mFopBiZgikBJa8YfFsFxdqEuFMBIpjJRgx7eiUoKXqPphoEaLHkdyI8668Vfts
Kra87sBj4k2REE2Xo91euwVJ2mOcab27WJ13xuvcpEU25LRqxrUPY6azdOYIzHNGFbNzvF5LIZon
Kgqe+ixYUvWDyjcCbpMmSOdZ47nYpcRd5Y46NbdaJIeuasFJtUYjm/focRGwKLUThCFVzn43N66g
OqwO/Ixo8SjH4rnLb6dkf1cYW9IAk6kfUvyAuDR/FzI0ALQ1er56Myt0h33pUfKnt9jsQ5qRi6T+
Tswljgt9fUXhz/VY0Xg8O1/PptA3yasRo5n7CGIwZPmtzTcRptm7hKMX1rHzZUQHE5TnzHEb4+9x
VHqb0f+HzoN3BFXSLUFV6P1ikjDa4wQYFhj5QLVfqBjkWM+hkf2r6MKyUQK5aTqiS2m2gHztJ5lu
fVgbwOTeOdRfauVe/8BPS1z+I2O0r5Ecs2azt2bH/3VbJHyGVwYja09+x5d/ddWbb72gavnGXOjL
Bk41bw1kL+a/h9vjmO4GIba8Mjbql8erP1Gi930zzOE6yct0IxL0MOyEWHeJx6oLJxsnfbj6gzN+
9WaOXptXc+Tclu1betMFaTXg5pfVSOSNi5zIzvm6JiMjBM94iMwBOjrMg8SLvdOUd8EQcQlDZUmp
MRK9iDOC1O1uo1h7vu6xwm63Ik8rmWEf1wxM8D2JJmPIS19bCETPIfV4kamjhT6NcWz11KME7u9e
8UltSQRGXo6ao0mQjgNlZSinp35Rr6RvEPJ1N38FV+g+fujCIZnHYRT2LbJIWwwygV0h9S+WJXxo
/NxDU0AYb3GiSWhRv0rzUfqcaW/tshImr0ZtU90+yOQLdBiiTMolwM/21aVnhC4586DjWT+kI2cQ
1hfEM6za8GAHlwN4EFgw7YIBYUrkVabhDmKDUFMNVE6aRVgh+/+FWu/X08BC3RPTjxN5+wPdo6co
npiLJNjtB9DgIt58VbwSZp0jMzqAVy5p1p2mor6FT/YV+OWd2xcW6ARWHDy3nShS/ihZzcN+4QQ3
xxIMHqNsr4y9DzH/qGPPI/MHy9l/RN0ewlYzF2u4aUWBI/eQF0DKHiB+g3Sjysmf/iqJmJpIusk4
aTp4erC07H42Ux9WzcGou1wXM8hGD/rBcoHY+6/CgB5RRsBy2isR9hyvYyjlSznrpGc4xOPO+X3R
N1jNu5ejVKpFJlLKsxalSbX3COA6djJuH/QvRYjCGKz7cmaObichmhx/5sbAkCJaxV8roXDJ7pOq
d6qtSxnn6j9etsip03q0ao4ephnHwKB8aw8WIRd52284ND16DcgbrOV05TtinSxa6DXwJk2y95An
Vz84Fwbjitom+kqceDLAO4+NK5EIbbZ2W4v2x7vRomWCn7u1Kgg8jNwCxrVU74UklXVH6cGT2z1Q
tKYdiEVT42LuLzDPUVeUoVwREOI1nQSWBi2iCOBaD21nqqW4z8sQpd6oVkmc1AmJs/zrEB7jRKHC
cCa7oONmti/+D+OJoIs1XX2HWyGijJwYMqGmF6KiIVYXrndXNa5V0WPKdu0Nf7+g627doBjHnHSI
kNMdAKVOaiT3iAoZzi7jiI4Z/31ZM4a5OMW26dtcm9l1JhA0RwkL1rzQ/SAmCy28WQJVDbkslqOc
W0pphTeND3chvVhF8ZoHqbnuJdaeaEjGa4bN0Zoc28mprgARp0oIGy8vPOBeLQ24k9gbNHGmSF+r
3nVWo2UXOZAzz4KVtqLm08jVCdn/WiKOW58kvwQB+dLTigY1ydYtnPPWPxBiykhbpOXYZKrr1RcC
AitW9QhwqK69Nr6BhGazlA9V9KcY008Xi8aDPn2QBGpumgv1bWp9QyVkSK7rCP2IDAvDaLD9IBZ5
L7SZXyLzVHPKihK8eIXPC3J4hVPNxplw/eQK6EVuoHaRrgwx9o8wyt9fK3NnQRUWXhw1saPnoE+m
ebe6nWBkWUqj/DwNJnhTI0w33W57yj2gBkBzEhmDs+CVsIz92DnbSUCbBCImsaA0hn2SXdlktALw
jnd+bCoxoQf5I+shsk3jsqEA9fe6GSrLFWw6bFJ+vJn37Xe2Futr1I6auNKz4OhTFxbnlgDCu4EF
jw2TuwLn8iQKDEunNfV5LkeRnn7F44KWPyHFX6P8XcoVZvOXkxZaIH44tSvh7LS8XfGHdwliINAZ
ZRF7jkm8bxXbgKTDoHyGcKAhW3Ssa0TylLQWNkhKABOhV46wZe/uM6yo5oyW0xUpH//07c6RMW3o
lLR6/psMkOkCSflCvBRntw2m8cMZuxbJ8kJErafCpDgw6J6/C2iDmjJXv+H107AoFQgeuXaSmXsP
yZQhnpcFOS80U4nLrBwafuGqhM443WKicnLCxhC07g7EWZcKNNVL1cTOBkbOPX1vCHJC/Mp3X/ED
1di0vlAXn3JOLNumsYq2RIa7d7Jw1kF2TZhDyaR5t7Gw1cDAs0C8o+BrN94g+YDKvggRoIg9VQNO
HKdFqy+CiFOKmjTfDkEfWdWdEMWxhZOwq3/JWFFW3J1TiiEVeQh8D+lYH/td/KL18cRT40uhGy3z
YuIStDFJlb9g70/0IL1wA0xYNkYFZVilOfA110ALUF/KN9B4b56thFCHAUQLz5liEhaFJCE7OdB9
SxJSqucB9IlPoiSF5HGabgF/DTQEp/XY+qU2UtbyUWiemtLhn23tePvpQa3mqdxs7ZOszpRZnUmv
WIpCKxGcoEWmmDC2H+woZc/h9PA97biFtbQOy7BmKK+altr94W5Apy6lemoJqSPk4LFsrMx24G3X
P6m1Zcq3QC2n5HQlCWHqI9D/VUv7dsTmtl9xXZID2BF72+UU7oLEvly7pxTSaTMutafWiOZhJVBl
+1m/WZSrsiTHUIJLZYMVhHjKn/DrzgNy5mpmFrJj6/4wZW1/jOvwMcMBX1mwgNEUN5KgdU0E5jrU
sS7LsTP+FO2JAP/MPgSsbKL4cqHIrP9839Axro2e9djXQrRsg+qDa7J+3fy5B1Fum4ZoAxRDxBli
yzNmkMhMwaOjjYMPJmF5+6jXt+Ou/uB7Q9EwvtPw6ih4WvVBKdqYeew/GUlJ9NVyilIiLUGZX04y
j3eE4KQXf79XWSzJ6H9UV43BIerpPtCqyn9PXEJQplr9UFYN6MRnrtFsBPsB8JOi77u21La1sd44
d4kMPQJoiXBsAOjrTwi8lPt55BazhAfLG46zJClBwt/srYPKjLSjnRGvjkizvVNUTr8LQl65Oj3h
p51x4DZgoGLN4ygLOHb2wruFyDcqTKXPI7plOdwRzqbLzFA9KdXiEK456T7yWBIODq/8R/2COCGD
h/HzuxFeTrNLLHDIncs6BIqNahjOEuA6/MfvLOTFOdTwjjELu00tbVpywZeelTP23RM4LpQ5ktWL
zsq8f0PgTDlu0aCS4lQla9UiTxQkg3RQvFI1Z/kvYf9psn4jDDrkV4Wa/2Zl9Gd4qSB6FEgttMnf
9oXEfMf4APwnMhM9bk1bOfpjCWvX9lTJ6lw8CITi67d1TPtxX/T/ZOq8sF7vyvnLHMhbycpJAJFp
3DTo7dOcmQAVgPKT57+uXVllyCx/ZW6V0RNIZ16RRZzYn3z+amkPQABvpzBnbHElSEMBIodOEJib
91/K9hKEJimUhWfzpoC5QP6uzi2r0h0Dt91FbY9JvtngYStRYK4ApIwwPybi4W9Yk4S/bUsAtEc2
M40OZ/NrgiaI78wwcf4WANu24z4Kcv6hMyZri2707CcIPJDoO7S4dvcENZmhBrCgpfiZKTdAOHq/
upQzkQsSjHzpsYkAi8IdDMM5oAaHzEXLMbxUF4GyttnNtSj5ImIkRJXMuEQpeDfIyaf0Ui1b4/6I
lQuWzemnWTl5IltcQvnqylthUozmC320bct0Tp1VwL7ZfO6yGeGyyXJMarMiItvQvClEDRBgDOUZ
uIDWd4+7t5iyBiKCX3E/MkgPMU0y7l3XZCHTcXU/vUqfAr4b+n1MBKJ42LmzEP6rnpJLJj5cViNr
c/kdeQ16HFs9TkU337rWLBvA9L1CKefsezkncdFBDySDc0Gw3+/scxwW+KwXHg08Rd4zWaacXoqd
+i+ng8ILGimXhQKRMTPeTYUPbOrotUVo9s7hD3CtKJ1JzHW1wNsQIObEtbonP3PoDopc2jBsDk4B
hGiDDo3M62vamaghuvTzIygOmXXVhl214lR22bnswp+yDZioz4x0Vk3ff2l5c1ftjpq4AsHNeeC8
uOWqqxUjnjJT93LNQ6U6TVLvlxshCKI170x+pd66DcU02uaUsuQjtF1og6TtrijeUuV5KtU/2tx4
532IbKeaXVMaRa555FcuIhJ0VpWoaWqpOEy9iBQtcncjRRHgzrBPyQPJkaUsrLau7mau/Mc8TlBw
8RkiCz+RPJ+9NX0tc4z/kRwGBMFb214Qdxe3IR4D6VnESCBv72ARygBdxxw+oOv1gu4i4y6AAMyX
S7BMacmIeHoV/3NHp5v6cjBqNGyCg9TdPc8N2JWl1lsALb2eYayrxQGjugCswoIKNmVm+kvz5zgi
M0agW78Fkt7/RqWYRddhQLkW4bwf6/Pq+P1pViB6GYiR+Oum80PxOCDj7OSyJrEOp3y/dExQvl7B
czrGXZ6POExqNDilcHSJwFTG7zCYd8uhcHc+9IqqGfG5ivQBH306dll6mfDBHZYCM/SjFGer6BPa
CI1dEIZOL4U6n1QzhR6pbGl3/I6y3uX4mp2Nmgp70/8o6ijfnr+B3gDxkYV3Uv/PwAqwTgqZkWek
2HxAKNTZbi3ADvrTcHGmEsB65Sds/8L7QNmf9UXit/mx5N+tu778hkarmn6tTrd5RT5I4dAdZljf
Pm41zi/MKsJzZFaClA2XN91ZgqhLFCTJdlNEHuNxsMvHajYzbCNF5vVY0nD13NYHi3NcP05kQBuj
lD/wQcY/fy+dtYverOTWpBdzXBVYINEecl875d2WNT0PJ61NKZsDH7DURAKfRH0vVz4/76Bk2Pou
cpiAcDOrqFZCUZlcNGicUAQFA6TSJhc32XuPRLbmoF+2T8wEtUnUT+j+Mlb2D+t3C6oZ9aCau4HC
joN6m8unjA2C7mnv/F3iOulO6UShm4UsF6c5P8WGrOyuTtWjtdfqXSQqhHgjaQULWhrguHxECq/T
7NteCEteYQ40YmmbS/clTD4B7BeDr45S1uHQcB9TLT0kGCea26Ss0RKM/OuS8BFZzWLfFGwK1gFx
eox8UjEe2OPDsr29iQsg51+jMXJ0MAJyPErBWEbGYgiRFPovDU2trFzEAuXQVzYAdDaMQzM5YRbh
D3W24CgS657EVa1nizPa6c03JCPWBPIIr0M5KCuT/7lF36o4M/Ye/Qi7GQUHQMIuWCKVk+pGO7Zj
vMAVAlnHLMhvwr+CjNymJp2jxdaa/KubF61DNtpB8U9HkbWG6ROe50ZZyU9s0GbZtftqfIr+FF0U
dCVzOjL/1wgyDs333vRkhW3fuO9him/1bCS/+ewuk+Bs47x/bsbJm0EEBfU1qkuo2PUtH45YTK9J
tvVV9muien4X5kSDarw4aqr9VIkM1/4IKQ9/ezw69mHAP6FfRmP/v6pJW4FcJnfAffP0UzWEB0nR
S17MWeg6iK6iYwC9ffMm5s9EAeMx4eXiirvNkYnuiRBIMHTEmdZ+M5G1nk5H3EmQTL0yuOAyccwn
fKNIIRPFMnxMddAoZSFqwXsSyJPkh+hqHPW2nKPwjUBH1M2ghWuZmrmjER4jJrTO2wmkiSB3oQD9
wOgLefAf9dmxd0fAum7El4JcoNzjZxHKBJoXP0IMkz/YLT/4WsVK426rlx5c6iW+jsNJpaZ1UX0d
pt7iIKlaR69fWdEIIRaLFB3ZO9of4inOlRNdEVrxHEzi7FDNWmvsXShwAyQebFDyji83a9FEwAl1
yO6ABisw3wNFZafCiumG6qarAv7QeehDDLAeL/VMK7yyKfkjhklmEZu5rUUdIE5rhHfoTDJkrHdp
A4Xh4oFPoheMZ/i8ieMWlMDhne/SCUwhzOx8IjIsrdtBzux9wnRs4WRwNqvBF+0L/utOnoTQKneG
oGBV22rMTcoaex0QVqyMuQKh7JKs7B4X574ZfUYNVNeYOaOyNU9AeOvtQ7s429bSid3op4ZN8r14
LJOs9jcuqmrghfJjrX2JANaSiEykxJ0qYHFWDp39atZIAGvAcv3zoiGxk1Xc6VbrbRUkcZteRDB7
BrBY6UmkKNntNPT2Hgp3VbYF8ElYpKdkg+WCNvI+qawMepUEi73zNXqgpVxjrdNoLipWOpeVb/M7
BJ1LlTYgtnRv0J163bZ2qVv2bG/17XwzhTtXiftBmhbEagPev3aIGtKP1HfF6dR3ZGmomRhQZs/t
vWNo7ZoIAjMdrwXNKrP4Kjayit4X0oda8/AGjObCUycu9/FiHijUrvt0Or8Bbf2pE73CzBVmXbJt
0rExbNtm9hysgzD6yP3Va6ZqTaQpl/uA7kpi+0oVnwNjGs1A1OlLi4j3k+YpNUdPGWCHjOBpsx95
pCofUoIWVVGoaihwei0NYPQ4xkCq+MOCKXiGVohIP50/guw7yFUHoUptukS9WTC7Cw0+6isW1GY/
/07vXbQyWURnSkRYhWeas5yVMv+tjxaY+NeCuMC+wtGw4fhGzW0Lhc6dJS0A8YbIS3a4G/cQpYfl
TuUuVLv4razIqcQX9pX+6H84E+QU1MMKAOGwVcYXNYKiSiSR7JICQT6tCoap0juSrEMiubgrzcwt
EtloaGBDDJ8wArV9iDeKabKhTcXqfdv3jUV35Y+qjgUB9rxF6TxwI/+c6KjXhnyo6224CMfo9+AR
lUSjkaPFs7Fek15VzX1/XTirdGFAC7gbuR4bOWzpaGzFcblbcHMeEcHyMo5E6jcW3QQj8ks5iT8c
9nBa99b4u5xB0uhGB+Al77RTJHv3r0ti/KIVd4fCizdegPChapnWbbqoJJVJpG53lA9j5IdnXK9u
3ptAh0+rP9PhOOYhCtCTvlyrWNQb+4gGZIoWeRwVRjgQgYy/eU1Es/Hk6Bd6yQ5x+Gvx1kSpiVN1
7RY9XOYgyYXDPpMn/FxwY9swgv14KgpF5qbyb1Va2/kv+vGg720tOe6Gr87FWZgWXCj9OAGsrZsC
tSHXFUu1D7mytNIOaodoor9r3tDouRibPRT5fGLHCsX2WwhbWRM0TXeKD16xQiigr3r5vXH77uQR
hAq/R9tsAyieIycsz6DLUzyw9vi14e0u6gPiZR866b8UmzQxnLn2ecuGrA+JUzL5m21jGbgJp9UV
tc+bnVDImS6pLdU7AYgziPteKCQdYch8fZxUV7iV1kpvSA2gV7ebacCvoZdW67Ot2IfU9F4WX00W
SaGM5RMnm27KtrVqJLARbUinQ2t7BGpM4mX0r60+BHPqbp9mF7hMce18EIbS/htGSLoIssNxYVPx
48I4MjuOz0rqOHPf5TzSKQ4S6bJPrxv2KvuL17bCLoHwic4H4zVzeDBVL2s+/Hyv5DawB8J+FM7Q
0OvBCDgVSJpznroUOO4f/DW8svCREk9nfwVPcDgv3VYyVRDfopIHdu47fuhMbWNL4I9IQv/EHJ96
0j+RNnID8gqvadRAZDxsSFfAKMusKqDM+viyXvYyGjguwBoMXsEHk8sB78KgU5tNpqL9pLyAIhPh
04uhRKSv8wJORYFqXF1HhktPDJLihWO3CwqvEXIK2KEs7q+h27kca7do0rQPScW2CWy/QnkAoIoT
n+V1J09J8eDMh520lWgUcS2kiP3VPnI/4KBvTLOhFdeqCi44SFHUO1o7LUDRUHRVASDyUxLapA6v
96FptAlAXdOILm8J2EwWqNGdU4t7SPGOZurkfRsEMZ0wBYw2U2gabT09pFVj+RS8LJVSyeCF4bV+
08XdhV/ynCQjDFNY/P6RNJeMKBU1G7kHucf4qqm6uhxJEEij7L5Tn3n0/32lFyDp1DXZPbF/X3Qw
VU2zOuzDD6GVGOqxzzSUvgPOZNJu9O3Y+ND3MiINaOZT3XS6FBjaCci/95YYXgY1BiyPQIQ5tFpT
68oHCnNhIXSPbFDNszgo7LxttW8eK1oNvrdJdNAI5ra9p0S07RLOWmXWbhVpGdy3nzyNdGtmiDsh
jthNLgM6MArbT9emokFbSLrPRdMP5I1btlFccJnZtSdKV6bYZR94Fxqv5DDDfXFn3a3rMZZVlmlG
UfnvmEzael5K8rTUr1MJ2Ev84UYgWSk322lf2gCYC0rZ+AlCB8C2BQSzMyR33CRFmyLNjYwxO7H7
mmmpzOsYr88gMcQdqW2KF3fxQxBwW0ORGrNIoUaah7t53EiyAcQCqwoNYSspKlrE37rrmc7z/H3y
guV3nqD6XGxe3YwqGimqi5cpeHrwDYh07lXJJnCVTqo+96/02cWefnplxAHrk21b1lzJnHl/rG+t
F0H/Qi0w7C0PzSqHZxTlgRmAevjOglCmcosZ1NrvUhU9R5OD9zNL4Mzyo6ikrhnqWDGYU2jMyIo+
0h3Am7tU7MjBvlE23WWc1k11yFzKcd0eBjz4Axks/PHlWNVUV5YrsappKXuknkNswO6WgcUTVXLP
JEQ2/UQdPW7Gf0FBk4uDeKh+z9cFgeAVs28ayo/WRihhEPf3KFjuKOuAZUOBIfg7A2musQkyJrUe
Zkk6wzI6WbtgF4R8rX4LdgyyIQT897zXXf2wI/GHPv5J9opZ8fKeqNieKywVUmk99y/3jpIY2Q3N
NASjJKFY6sTd/mfxUDgXhObZsDvVkEgu5tcGF4Ew6zB8PO1qRQmsI2460dnl75uBIRcl1KDLeXim
9JHi/F7nGiQK+V3XGUT7sK23AP9HG4uNEaXa8f8hZnzjGkjtPjh5tAjEFblMCMiVk1pOe/yQo0PA
jHrJ045IqskYAFXW+bupY5JU0yEtIBGFqD6SggyEzXkBKu39DP+9FrSLJUHeUWcvLx/0Ae3Td+kQ
8S4F2hQOwnXChiY6P72S3XXp065O02Ldex3Z+l+qbuTn1U0rA4KCgcrKOZ+yBMB9vsrGNEVvvwf9
n3P+Xa/BgCZpSG5tjbGO+VHLFSTLYGWFUWlU9gti5Ml1jGbfIccsIh+rwBgE9dGX3aRMIzXzOCSg
/YFmycWHxmfE6/+RMOLyrsu71D2wMy8aQgAhpoVTgLZQzkT1do78KdSG9X+YTR9kgI53sgVmfEEp
SkJofUKokT3fK4HhUmygVCl/NpoWfw0soKpdLydgNe1kQEcZ49cwnqVcG3VMAIRHFcr4dvhWMSYf
uLu/UQIWMK6WdpwqGxG5mKQ93etv8FFK3tsGgT44aimgosiAP5pwY0+KBWx+vpeeVRwM0nSdvXZI
Dt13BDJdldNjSrmB4av3mzOtB1b5PmNyQUWzXacXqCYR3EGI6N/5IbL4MHXuX6Rdzm0OBQBS5nDj
ouOUFdCY2V+RC+AR5CDo3+oCQKdOULU4xcKdhDgQ4cJ85hr7/xf19nJASqwGCepVmL1fCFmBFWTx
pale+Ucgb6H1RXKJbLJcIw6itzX9pxEvTDbNJL8yWH+GlSJ7p4LsYhBdybW+zf01nNrLNsbB3CtU
2gQqZDoAWMfAP/4DsY0r9G6TZ0TF4IHyFS/A90aAfXks6UbRx/Yc5SCjgIjv03tD1LccMVPo5sfw
8QXapV1C7vQAhJXqArdZtzD4y0Ga9bBc/YmHAWkdvUxm5sSgqBQznT4qUdlm4hREX3Mc/eJmJ/99
pI+KOtGEeRdH0wKLFWpl4rF3axS0vquYRulqWy86cdkeXi/mTBYftLlmnHfeb2hSEWCU2/Kyrpim
2RsLPNFh2kdgUM0rh/WXlr7swP1aY6r+T6jGr7lYAKaHyW+jTNUkxtdXpmFDh7prc+FgDv9L8JDw
hy770AqS5tvMjv2p+4yegf/5fk8rM+IPll0lvIyLI6/FJ5+aTbBjGXexwjOPELCFQVpM9YbC6EFz
hbz5x4P5ffsC/bc2nkiTDKfkp8L0WWl/chXt0tjI5T1dyxibw7fRwKoqDP/Cvv5+z1moPpGMWl3k
CKL/shtzDlUDkqbbBKL56hRjjCrL4suGzXYJaplXXTCrqfooWLW0JbY0HBWDNeOc3FcIqvhrB3WI
CsAefgd6HOGrH+s4hNj6MWX3mgTMtxbW95FszPjQgtbOLQUX0P+6zyjBKlOtHDZwH/yFYrovKnlA
+rnIE4CM8ptVPeBhL9vs10hAb8+XlYr0R0K9rPAVgRGCaIi+cgj0TAsl1iyWZvbC8lx1LaJrv01S
lJVzTftUjpfctpADy0b8b6WnMHZz8/cfVVAvqMHEH+ZRbvYDEu3+xwE6XE2xMXSUrwS+xpEs1UOy
EpK0kWr6yQDxu4zghfF5pcyCGYYgmXekYqrpehBbWpzbchak27J5ZA1WihQ74Is8EzSGHT56t9pI
oFMPQeZkYRv5KJl0T/ed8V5GqxZMRf/fHOYVNTNDqUDxxD/JF4PpPcZAkWW0miCLTJRIDuxpEt1B
X3wXGzkdpyA6SYMKvijsaSbYqDbU7eJHg+HjZueMevUcQ7OPXfdCLVLw5NH9lcxt69DZEiLf7u8A
tfsjjYifP9CUA211GXbsGSghR1QxKahZo04cld2UcNgZ6VKafiU22MWaIZFi2tokvX9/RNxFc/DN
Wnu9HbGZjdDAP4odbNuL1gRlfC5fEel3imMjJnjUbJ8rdTJKW4WLB1OHHdl36wJ+xw1sX3Ye3YT2
KyHoouszoahUTaQ7ufRe8XNlLIloz3ldhvlhPqLXbhkJv1iPvJY1km16CTptUPXdoqxBEUBcZYDw
IdHza3QjVrR2LweaKnL7tdcua81GKrbLnDtmdlY8WtqeX7oZW9T9X4jarKCBgE8Sv7o13UU2Y6+u
it8E/68oeLsucxDochSyqNn6qyjuljU+Vl6KJVCmfUdABhglpPztf9jJKtujcu5Ml6anC/DgM/1f
mo7AAJr2z0ApIL+MtXBYizqAJ5DFnKG4Z+h0fIPIaPwQ8jqEaJV+3NMZb2+N9I8lDAPZbAGhD5wc
djRCHgR2VR9jN42wMdnJqHF0mfodoIOzDkf6g5Q0OS9ioWwcMjNHBwGahKmUR8BWDphNHgUfmcbq
h6pLAu+axRKDZ8B7iG2XRZ+tvzmk05SdM1SC1Rskv1Sozi/3uH22PSXYBhC7qnWoZUwTa9Yz4sVY
BrEZXJ9U7E3+wL1AxyDz13KN6hqwLmYuj9oR2d1EMxFvSxyhKput9DgiS3OAkc3L8zJD0drpnBRB
D67ot7pUwU5aleU8d1fOUvVcA4Wf4gDDlqTuAOb/Ti2cXFP0W8ujLcDdCsFSXgBdKm3ZiYXVaKrv
jiBDx0DqW1k0pQQQNfvfEjm7tzkojgabv3RFmpjZxvXVKUucBtU72MiNe2kG9YFi8DcTavsrnDYZ
X0TF1YxJOHgctIYJqKaHSqIMBIxNO1SbMDOXArdbmeqv5XZX8EUcFDCUO3SQDS7JTzo9H/on6NWW
L2qE8YhJRhDwSJBE+M2H3QLr8Hi3VJMXmo8F9aBQmLGW5Yk2IRsPsMT/4qw9XXSGx+rc/iOShJVZ
wlBuNXXLRl5mRGFNTxd/8LQxaSyDu8wrwUlfwWV0INlWzz8TvEWAeOlO4LjZx0Jr5fQaltyOl02g
oAT3bzTAgw39luOV77VAxwYy/4HdsBVpdwLZl2r/q2g6gaokSUIBpXNUGDiGLCO8luBEMZwaglYE
kY+GfBQ6GaXX86g10NBQvcpi8s8xc4sdmkVNbeiZ2KmystVoRnhEVeAGoVNfz/axf1c6x0N0hIJj
AH8vPgd+HsOEq0iVa1u2gK9FnZOuOk9U1PlkcfTmjTCfAy4dx6e/rXB5X+i3CVcHSXx3Rglff1SX
o2C5ntqiNxfz3MRr2Ezbsw2XuaIH+gIvwZ4PT/w7QHMflEORFHCEGEp8EPrFighisuJ2SiZAfJ4C
xPiw2MNqYvYkHuJqVAWILUCeb3UQhQyTsq1JRiuP3cMApSwx6l9BnPcu+1/maUoyMijFry+p3t2H
a1IRT95T0/1A2idRpGwNlFF3heBVkkV7w+lQueNAtR1lzQzVaYXLDJCQabbfIRrZqBBpchKczuI/
vmH0f37Uej6seBfDwTNr/MiFabeWxmq6fPCdgigO+aHoM8a41QHGnvwTGB+toUqbklFsOBePcRCz
jNDbhAvfbWZrGgfmjJz6P3jy5w3P56ppFTG5sOfOIzJ5CLk3oBBl87mX+gj4TsRONIMTrrLckH6D
XINpFXAQQXb5O7+tbFN2gmpAd3M23Ro0hDhDAXFiN8ZwC2HRjtuwmP8Q4rOvggBzChOY/VLJlkcJ
a4jzBXwrbv5FXNVgDbOOagdT8H5VwzCgAi/JKDijWRlk28rw10r0sYUgS0yMZFqdTSpoq9vdziby
BLGRPfGNVzeo+oojIYDvW7FVWvc9rkm/qftukHZUnGFZuXaesm0r2cQGkYCBUGzrc81JX4buwwyN
387KXQ4bPMc1fp6UgK0+KKd5hhd+lssgvkFadlCEfX0TqZrCSKQpBBewTVvbFY07L+wL232Tt8+Y
pAV5VNlIkaT8/mDtSVWPTcrKJEO1y82o3gKl9lWG0SqRee9UcHXa4I5UjujYwikENj4YmaXWA6zh
I0YssgH+sqXfbscviZIOj1ibclY4qnuYpyyGlRA4t4/TsjpKg3rqkJvyylD74mlVRmngW8dFV8dd
2ductfL+TZHhg+rOZ+dJhZHDw8C3unjfM+TvBxoIrXTwQsoCnR6T8hs7Uys6IY+xVd5ZH6ygsaMQ
SA3i6oI/STxT8cQ4uMwZUoOkJ94phcrQ9Tja4PBFx1Aq/ReNHVMjQaR6QNVgfeecOZEbkvs3tdGJ
jsOJCjCqKr+8KxrHliJIRbx3I4bxD3ScApFlWwIqOfEovgvSREgW5EobDpIlpaTBSJV5obmjrCdg
jUV8yvsUmQOEXWv/GxPHNxqLdeQlbmPw+6WTCOtk/4hl9TkvWFl6SAj66AWAGieSpBEVp7I/Zayk
Q1Eq6S11u46INWU8M2Feyj66d8QMuOTGdRJ1l0O9X3v8g4PQOQBCbnQ/UTcFb4tCCObicpBT4Iza
c8RtScnYgv5j4WdqQNZXTQohn6vZ0Bp4SZF3K48+EWqP1gYumK/4lt0/c5jFmQURZFiVJnKTyyQE
Q1+rdaFire6x2R6649yYwA6hteZqpOv2g2WZMjUP4g4r4I7QWnifF+jRQuxKVpcImU5NYPKA1RoF
Ru5eUHWhrwcmpDV8SC1jhMfpo9yLuPSRKnXElE+GHXRZ7B9qlZsUJO0aN3OIyLuyB1kMYUlk4/Ms
5PNO5sk6K1Sh1AxBy3v8OlPLZagOu+QcQo47mq7NhMOV+TZg0NHPao7bNvZ3maQU6kCZgkUQusu/
x5oxG9jsvdz6th2ouEQWzX4sRYwyGYsdo4kc+qy5iMbPQT+3sNCmC89UIPLD/Oa2qKw/GFEfbQX+
EcPP27mgyeJCYDQBLQM1+wRADGwKdKUWGbODpM/tlykzAdm+Q9clwVk4aB/pN5o7jsU5PHRISnU6
5Pxu8WQut3rEpRRINHO5KDdkvmWOPOq3Rn6/Lba4jih96k8008QmOOTeQpsM23j0jS0fVP6pmJhe
oyGEvqNh3ysiJkWZPVoCHS24P1TdDAPJVvw6wpRhMEVk1uTPx0LyqSyeSf4L3pEqMFXuoIvfwr+q
5UQjB/FinHI4wy68w9gkWIWbLTDk/Q6tfE7FlXvMP+zJBrhqk69f5LyZ1iQqDAE7GsbA6qumpbeM
FVXHRz6P6f+SHT9Hktic5sYdw7JCrCfLHZ7FWXQO3mXca4ZeuhIK+OaoB+pLA7tqveLsNiQktxKC
OToqjE7tylI/eTtHUX2ilYtJhqYCxRuSswawc4CiaBCSDDAsofpzwkpNhIsmug2i1I9qLv63BSlb
0fsfSb8hVArqY3Q9x77WZJ4GyqAEw0fywvauT9T72JzNVuBMR3KLWVHFHxtNZGZHvlWX0+9yD1RF
QFLWtulX8K/pxjPavfv3IYYigIT6vzdPblNP0UvjOrnJI0g6ViLNYRaQK2PNwE3yhNGg6tJtmr+U
MKkpVJzvI77mVtMvG4AWGfMtA9nfVb2Rncz9aaDXkw7AkWz3MRgNoeyYzN/kPTHsE0hOYkUnS2V7
+cekBQ1Pim5XXWFTvqy2AHnrqGi6+BBLK36CSpjJF1kxqyubfw0N8G3+n8vu8hFoViRGB8Q/4mJn
2j4okI0ZDSxJkAEqqn8w5UtTvstqK4HHr0GKatI1mUL/aCkAPxGRUQEY6T/tLgrytzhu6w4Hvf4J
9+qkRt/x9OKxGK+KAhw2wEacObo6e497birFU5IHwX2lzhlqBH99e339MnPvqg/sWG5+SdYRTq+B
eajF1lOoXmbWi0aAFhuUFeCpeDf6fzjJeWvPYqYjXi2HyzI7UO5n6uauL4Wby68tFblwmrKqtgQh
8uLkgPZBx9afveejSJgnXt/YxFc3liHfV002y701/tcjV6baodHPR1oFbWnqbBZeFuMkvPRk7Mme
Uw8JlVLwOYQWoRha2lkITjFLhhNx11IM4y0uIqypTVoptKnsqemsLXaqqd3oPC17objlFVWeKTFG
qzCcFNokpRAAH/xKlyoMPLyY7CBrXUdggfA5iFuz6OMY2KhJMjn5r+aGHQnPwjrm9iJ8aVqM77zA
lQhZZUBYoz221gJC3TizhRnRcw3MQErStirM4ABiCqOTSwWSLBrz4gGwRFbuaaVuCGQW9d5cbu5G
iIoqF0ZumuPEGCIAPq8GYWetTe3aZ/bqXYyhV25nry9k5pMHFPZYA2uc0hIGMVlSUMLHb4RS1c6z
Hg6yevF2eTNR8hzf2FP8BgyavVD4B/uhC3eKfRvwHrOT3xRPXnt2BdCT41jJ5RO4tgzO9X3uAoP3
F/9OO4MsMq87IPj/iKV5KiwlgDSg/oPAK+OuLPSqu+7+5D6YmHtx8aKv8GNC1gyYCCl2fDwozrdE
bgvypYm+OHptCUsDAt4oe+ywJrOYBwL5J8ZVVkT6AiezO4WuzxuJa/Jk3ithsKqeQAwXEiQrz79S
sDFDsUuXifdASeZyMcUNUjhgzSrayeSg5epn/vDZoHBpL+0GEBNpaxzptlJlpDprZZmkua6lFT0s
L6fXQDkZ47sbFtDHn5PTg2ny+3h7FVRqpj+y6a6p+ud+J7ZQxOw3/dV5uG4OKe6Id73SGfs9ZT6y
IThgluYTXld3BVvD2s8D5d5cL8sG0h5jCVup59lHkwKHTiHPQqKynDY2VXjVpp0xkkWbrj+T3BPo
WQ5vQ8Au6cfqX4nXnYOhrIxkFPlJEcmwzxyjbs7RF5tY85oqKS/AWhSAoyPrxyxJKG3r8TKaUQ7a
aBLQr//2SG3JOL4BbrPPtrX8JNeJ+N7oZ/8ftkcaJMY6SqJ7z/MPMF6sZxHs31mTI2PqbfKdQ2wy
TX9+IlqzdYhplzPBks3CySMRS+RVZUhQU+uxtOHJSKEHCoK4qGNQ386EYZ6MeWpBCy8NTrIMr2f6
2lO0L4C17dywq/x1Lha5EX/3kTX/CX6Su1znxY6hJTz/vZc5Q7hctSA8DuTMT57ShIowJVyhd+DP
mmu88NnB9VVICkgMzWLMrB1ix3WQGsQIDhcMv7iHMsjuCtyRjTxERV8ISKehPgmZOjkbs/VclUZI
lNgArHtiYU98fj8haJ3yO71uuo7mmuCljI7pJLm3kTHsvNMJcCa8A80ZnCEEulaGegLxv4347I+O
wd4S+w4mYV5/Eg3bWiflPLQfmbAYmRZOCQgihK0v4QrSnCEjOizko5tvtakqXUgaqABgSVxa4CE7
OfnQc9U9yrOdyOhMGugznH5nmC9tzZolD/ZsVu4cF3IJye5bQtAAPtxDDw5Y2K7GVhBkKnbjBfdC
1AhtFadBmBkyKuQiLQg8rvlLMDjLAaGXytqwTT1ZCcszjBGUatU9mBaG+tFLvDb1t8rv2VrECjSB
2w53jcZuRxlXDNKpvPN+VhtC69/kZUyJSdWallyTa3KMRQVeNbCvwFde/BtwjfNGw8mOBSGEGWrE
OqBJ+3gjo8fmAPi5eSReUhIjELTwEdslrEMW6KONbruJkMs7wCl6tvhw152TP9KZUuDGPlTxePgI
knR67OG2vjrnMJmRrXlLE4MYwP2nssRN/CSs4c279gNsHt5VIfLXzHQ9NxeTgaPXxcZlzZu3sBE5
784ShCTO/zbc7EWvXKL8dbkrJI0R1KJW4oEpspd2ys9iZ9R/JYMgEnLxtNxuuiTS4Hho6Mw8yKff
9j7zfU+plSBzkknP9Uh8AdPXUkNhOYMykdKhsGQcK9Jug7CjwKxN1EEPwgqLDJN8Cr4JPoLdWFCG
HOCpWEO1Lp2Cm76EMzJfL7sUxvmMn7eXSwHRRa1f/WBpqlMbArRLpQAyz5FGcVs3eQENW58EayLj
ADGDGtAVkYhiIUiWWAvr8qbu0DEZsugdR/KtCt3Q1LOrBzTHXy+ZmquicESTIrUyF1/AfB2wfKrN
NEXVdjbZ4gJosUhMOBW6+A66sH6ZPotVBDC/gvmnODki81RRbkv0c46IV7MUGw3duTmEKiyINMLu
We000l2c28+FsVRCDERGLRP20gGOiAO9myVZt/GLVs+jE//Mbq9wNDrlQ81BxcPtLU3PWg6OCzZT
NaalzQk4YlwTKmL90U6OgUpBhkfiw85YxzPub3P5aNdjF5hVoioGyVhMqFlgkfqnkSM2wgA/UNiT
DxMc2elYLNF0DYIsgzFeIjZuGMZuA439cI3U9xsA1sB0TkqvEdeTNBcY8r+EXwfv8wT4f5W36uyN
QJ3CSMYUd+I38R5p0ApdFHoc/Ms89vRi9Rgj/ig9slHsPbxzLVEh0GgTv+iVN5tJ/WH9SjCmp2OE
QHF5PQQypJ5G+PzCOPnkg3bRC+5J8QwKSuj0tNlyPfFlbJfaRqJVIHToXlZoKsNJmnfsHitC4rXi
SOZQcqYfT3celcZeqY2mENAGi6Nrgt8ztqX19KzENXB/HCwk5HvKBGhP0OkcVltQ8kZynzn83ylJ
PyUOUgLOtxC8ofEdwnC/OUsi2uwlBk0GPrKLtryvoKEKBIqQ7zU30EhLJ1f7hco/hK1e8YIjMunG
MP0qTWUE2wtQRWT3xC1C7u5Gc29o2yZXbvpVqrMzxCxNxwBzCTGzvwYI8zrNT1oSXGOgXY4fQQcU
WGXRl7Q7EFDer+xnbtz2JCtGivSjCQjHjnQUWkU+34N9BVdpIDmCKvFjzkuGJWQFGdjVI8XCBy4f
7RobpPxLfhDbpIqji2uFgRMKcXJG09xcWnx/ZrBLr38z8mhGpzw4t5013Ycw+oWmP8Xk1kIRED10
iqKog/8asbyDHPHkn+sUH4icVs/GkxxI9TgdBO+tyGxMQ0Sxr09/oz0WLHLFc47w0a5Ai/pWsE6O
w+79b7XVBc7R6WJCuaKeyAhDk/SWbWQ5NRUuXq0xI2oN1QjdUPvFT17NhpT1kADQR08u2jbphfKN
Ig70EPTLmVg8a6IrIrESYkSqvGDmEJkQJxOb2NjRyUIeFlRRgv4R+aowe6LPkijNTaOIXyfE0ULs
Aj2cSCQQHE7uyOs2qPNKKV//ibmAhUiO2vwAnrWZYJR+FOq9iUscsSRD+cuaxKuyvIvsj11Z2BQS
ANm8mxM2qADmVvlGpLkfni/uIqFT3B85JQxPJZGQngHJv+RIGTst/9r41dteYRuhhR82T+HzwSoP
6fyoH05V/dFpVRunSB3khBa/gceJ07jKnMM5sBJKApR9tK6MAKWbKs1Yyonkvqx4vxtOyLIc4QxQ
uxy+SuKHZgdV+JuEwUTxtyc9LCrYtcD4Y4yGQ46STNXWfVjB31OBTWOuM4sJgubBI/+IKJf6kNA8
buuQOeL+VD7qFyf5NculizU4CmxzDQ7XXj1qlj5KLeUXDMIM13JwO8ztdEzCs4rhJpx1hB+9xEtr
6OTk0fwf8OyDZBzIYsLlBYW8p2RY2Palwdq1lwmVvi64q8UdXL+/wZ3vAUqxxhNFice8sVjSNoNm
E1+wzTzmed5X6dKmcbnMDY8X8hTquJcsbTUz3GxvdNfHCp7r6+SuBm3X7HsdApO/lnWCTFPGjdLX
kXeTdnD7GYcLQzmx+mhJhK/Jq+kh9KJl7yHgAVwl7jEVK/Q8DaLbGHjpxnbykivTk4wYE1Y1MEwZ
zBs/b7p4ynwnQpu1/96u6b/IpqZTHRpPdky5YjH3Yocmpib4/J9E/5pRF0ESa+ofpvZvhgjt39jQ
Ae1XzJrOtSawLRPIlCEfwoemHsrwbaQJZxCTStLynj1Sgi/dMmIsBGsaBOvz97Fz4rKaV/dmYsPx
zpJd6srOmH4rgSkZNhhk5ezhr+jBzKa6NVe3KRcJy7+O24dqceGM5vUdkLaEJTrFv0xPQnMIfzsH
vIcrHe41rMtu+SyKcZPc2q5QJjJ047ZYGcO9Qz2wfg7lYH3gzBVI8U/BUloKhlD8/yKfit657Gu4
aoMDS/faa90ap3OnMh5thVYR7MayM3vQZLEfk0uUa4MePh2tfS0UbLXkarslcEE0W9sp/CXxP5uH
7Xn3vMznZFitqCDiKANm1LCuddEfI2prYV9WxLiI3ldmxr93+Tm2nMLWfSLqopOsA15AZwRsxzGm
TEUcERVIGf/FuXvMUdFjBrf3Kiz3wt90IDUuGrJPWbN22DoEJ239DzzJhyOuVRh26kpK+quWvBE3
UGStgvxEHOFnYHP3dQLHeKxYM1eY8U8WyjMQJF9o4iHef2SrmX575hp97/MtM8OWgzXZ4b/KkDNt
v8yy845coOVksBginucujeQud2mUdpPckpVygZmjcEYnX6o+T+LTdHKGJzzbmer0TOID9En9+glp
386Dxn2UIgYx725hxUftFRCna5kpf7uFXCpuMzbK6zNKFNjGE8l5CPN9CbsmxsvV5jF7Y1it0j29
Is83IKjcxS0P/fVH3CHvzi2sL3CqT6OM/dp6S1FPA6rI3zehbtUvf3n15oNgaP2BeAo2ql6iiuzZ
6xs6WyfDIMML8mmAUI39IKpX2NyhTiMgZjHV28lqUf2ihgmF1kPpt8WklJtOYYvTdY33pnkrKHMr
KVgn7Cpz0oj8mR8Rr64wU4/6bzvPtuaeSlX4MXptFOWHWI4angfLs+r328JjtVH4a2ol1r2Blwi6
LN4UDOinSOUrqu2SYhSnyHTOd+Epe8ieIOl27QXig0w3qWg+aEDep22HtnErKf6t4Urmo80q1dta
asOhdgegs4omdMSJFTJyLMpIkKAhXOkW08pQgE86Z1CCcbiBMvWxzFlKR2OPDWkqVFp/uVAKATDu
JyUKqn/6kURXiPy0VqMWOgSFiKu1BtlXfpFuz32idv6+ObTLGS918NvvtokRNUvnxNjmJ3ej3lzS
UxSprvh6oBP4kER7FCbelJhJGIyEILoYMA7oXtM9XBIjS2vAvPUFinSzBqSCzt+RH0q5bKytEzqq
GjD6o5/VSTgf0u5jdT4Kln7Pyj6WEvYoVNl2WkKQ0ZXaol6nDE1s8FyxbwOHBoRWYt4SXDBSZk7v
QIO/abGvhhdzOz2PGPeBxONPwco4a58ifJ3ZYBJIRDowv5EGsmArlJ7u/9wSRXPUfYp44QNIOpOd
4m0lSXDo1fentQ5DbZUVj1cH7zEgIN191bLmWfFywq0xncyE6FSl3DBRVtzVzNJmYs1BQb76WryN
bzOV5BK95c9nkeKFAVnnSGLijEM7yhr4nOQwrut7p5/+w7o3tBRv7ZA6lqtmf22a27nOSwsdNJoO
hNpOhOvrh2I4hdDVXCKnJE7wkLw/Sqjof7ora3HDF9/ivdx6DKsFK3JHrw8juyYSBM1lG90Uo+Gp
qEC/xcgPvmC0BkoHnEyHsRUvzNZ5HTBThHqzPQy4m862uYT0KBZMR4zzzb5TXS/euJ9AAjGwW2gL
6A0VddACJMExICBkbzZiWx/vNNjOPrPNyodeMJVxoJfQqCSAHS16bbb/xyAScfj4/IiFTUecW7W4
tR3Bql0daj63JxUCuoqMYH9xzbrsNqPmePTFvOwsZ5YfkkG7/V3ZjdfZiivI4l/VgdvhLNPjmv1E
MHEXKlnea9nMNd/JjhG4Ls8ggS/zHrrRX/QuIIdowterZlOhqSVx4XEBFO4/hfaGZOb3oQidn7VP
crk5iTrcwa06q3yzfkoqOQ5VFD0XCxMh30iZ09TxN+LWRKSNOJ5QpgQPqyKtfuoOoj379que0B6m
uAEmG0ve49B8hnHdWp2Ixl8iYK+sGDmEpUbKt+8PsCSiOts79aVbOxRc0g9SJdgAI1UubJDsxp/5
vUJsTaIWIVEDob4vrGAZ18KUPfpZKmFBBw/L8GcpnM24ZQxeeK8YseU66Kot9GUijTa4vQp07yTV
jp36qcbopGMtoCRKBhXYL0uR1oWu00YG7Ibob3HHucxjsfXwTR0Vnua7IRhu9W0cmVC3qZ6WSDNt
d4sHnOgRbJsA4bue48IbaYvioAlJArsdOPo8vBUxyyEljGh3sDpV5gR+l0+7ohBjXDB7ZG+V5tts
uCQ6HnwJDSezK9eLd3yzd41C1otwvO+0BSBSoh08MJGXWTDrP1RlVH7f/ytqYMpLuw+Z5cdIq6ZB
Yj+8YHrCgil5mWfMmN7hLCYvI28zBH9mP786br0kpwsI4xIPhLtge0VtPzPmC/eQbjw/xlsxOsC7
Hj3f9b9qI4u0NB5kFtHPOUovw43fehTQNWdZ5WNZjjJKnY17NJ4Eew4JGOPEvvvX1YEsJYqYa8YW
gfc1QJWH1nRAg2wY+jZvXvmqUGz19jHYdtaQogIf9ZHkXIIOKEhCKnSHxpbRUhG4Dc775rvUokn8
HR4DmQtiO4VjvAtueJiJZGC0exOrBi8LxBSjFsLNeDoFypQhEIDZPKAKoB0fbNZVm5FW5F6OH8O0
Yn8BsELNqzVQneWZGbJ0MB4lDjPlQOzX9ofWGkmG2U9MIm3ueBbS84Zs9by2B4f2C4DNqLFCbkEz
rufumbyuG1OUN/sCXDYD4kCSyy+wqDtt8IMz+7U2VIO+rD4UmHUB4bg3ZmJw3J5rIZpzHVXAURnE
a/3lDXrom99uWYqGRXiN+puMzAm55dV57CCuzAWu1Fo5g79MBSX3/lSFvYV3TD0mplnEfz1gjcOI
AFY30W+6tefPwtesdfJYzjhfK0sUanw9k8EqsZACeRe6vvx4B/Ym9jsOjLkL0lOkRlIZlprEPbvf
TqF0xXoSMjrnSrdYB+ZGHHmtaH2rN2wQYlx/GYoF7fBWP/AY4QUeDA7it+Wh2J6Nu4sJkMgCjJ00
DZOIhn/9I7GnhkjwKo3kZ3nA6HbXD+PSUBffYW7Lipl7YimwGEANM428E2MB9odadyO3oRN+1zg1
a6ylH0cKW3qdWRHhfRnPRYAVd9YrUuFQW22fY+fUQ5A+3SGyU5D+wofOTvwTo7RqqVocQwV41g2R
VRjFVYPOb9EH/cUHh6/vIhCc5iVz+FOPCl2Uu8liWt3JB58JgZZqRbe9O2Yc/+R5cKEQXkKWz6oB
MqrimqfA5f3SLMjX07GFQbvUyAYDH8gnQDFAs39QMSLxehu2Z8LuaP9eVzNH+CrsjdwzepZcSvTL
q8+gSKg+1xFCUzShK8+lKOiG6rlRWPFGVu65JWrjoo/cncda+rJvVDZsKMtLfpopciQxPCALb7fw
O/WUVxoQUnMKUfKaDjVm8rSM15XAvkHbXL385kcZD3GIlEhUXmXbBbuLXo4s7/5AL+N9ZmI63f4J
98ocAI7yAJmLQA49HyIwyaPZkiw7GZSYGrZvXan0BjJZJDrcOGFsO1rSNNd8miQ8DvyFfU8INxOG
ydy0nLr78HIdrkjKXC0fBrjerf0ccO17c+O2BwojFr4dnoptlvwW+rBC9xg8Be5UPrs0zaPL+OVK
zy9P94xvVhGT8mgi71tQPMYN25uIq0LsdedbSMjCqN368yBUgkqdKBm19c7w0qbjSZT+kAgTl1bv
Q2RvQ6Sc0lwVar8VFAqLX0Q+gu6N+2LvH8BQl7zmX5As5hX3eb3PVj0gtOZpx0SGUmnfXcEtIfKw
Y54lJ+V3WoT9GyMuh33KcQascZIOjWaLg3Ai8KI0qAMzILc2a5IlMFWpZ9JANKl52E3k/dzq3BmB
6XzOypG0muIRUx+yKCs66g760pcPWRZGZmUlBoLu4LnWQSjRyRG8pxCj/87Kr+phgIrKRSCKyTFT
oduUFIBsimBMtXhuxcgGHn5IooP/XSHVLTS4/jx+v29YTRpn6gyPfY1XSWMlGOq9bKJgOYrv9ne9
lF48Z8WxWscJyFqp7o1sQ1iK2Sb1qwGaLKSOloI0RlHRO+ceLmY3v0TehkfUQvrgjypyQ2SJQnVU
3yujK0wVVOHAqHUGDIBl0ok6sAHM6uGRP149kFgqCUwJJXNCnZ1dYD2wizvSFHlPrnAMeAfan6H7
alRlm8L5Y7bA4Xxz5ImtqTg1dQvKkLUYErhC5G44OsJrTN5VAHS3r5owAt8kU3GvyUKs5CbiB/Dc
KOHOfrTNaGonX8op1Rcz3ePobhx48Adp0Oshmu99H3q8L329hMs17xykYlHUbSKyrmC18JRoHKv9
SJjG9u28PHDG1S1os+6F1RqOOsvhJsy1veS9r5+rb94NyMmNbQEUS6mY70J+FWXqYrq6bgithpCh
wj09O+F2ovwhhUG40D+fY/rQdO+Fv6EkFsn+++tndBoB/YIQ736nOpRo/SVSxlEzEru1ko9xaAoK
ndxO6p4dxsP8paaM1tMzFuhVkVpckW2CMPxvwBILYTqADvIuvZ33pmleJk3BkXRmx1IYVoQmY5OV
mKJIfub/h0C+R8TiHv0VR+1+lur9r+hD+NOy7jLx5N/o1EUhU/H8A4a8jhLXwj08uRhAzeijpELB
2fJwgQvSDFIg6Lsf+G/ihcqm/JFriLZtOf2SIijl1YIQMX3du5VpRCLEUoxMToyCIByy17qPoGac
7nOCY8Dr+xQBwqTQbOkx3Haeu8/CpbYRsnsr8H5LRUR0nN6INvKw5kdx9ezngMkeBOVP7HUy1wpU
qUsZj7Bxa6H/bV78OYtdse38CcfRRlooK3y6O39yBMvBTp5Jl0STz9NYtK3K5jAiNt1OyzAbfJLr
J5C8CYm/o9K+/R0IYFnkTuVDPZf43CddsGPd1bB7uBzlctChTgqOsnn7nnKR+dCZ3RRpO19u4fbt
I7isHq60M7mX2ANNQORRZ3IOxdPYs/UJDMv2CxqpJqjA5bqzsweVrqa3iVzkgQOSnpYn6pxRK1qf
PK+s4rXX20cmdPi9U/4/pogM/6EokPtVF+ShEIsgWOvG7/oDXkxpc18BN38uDme3L8cPXqhqASnB
VNzW5w3vUGTMK53km39HfV8ZHip2IWHOA35h9/D6aJHUD4PEvWU+OdtB4oIZh3yGkhfEqN0r4L2T
e3k4r9RTja6QKnANtSRUvspUINzAvBKcqCnumek7A+gq1HhDAwzsdBZMQhCSbXfihu2LfN3Caz7B
Qgcgm53Xsqpz6L/mU4RJv61kD6pA0YmusUxgYXC0JEeJbHCcmLNbq8vTFvFdjn1r/4g7mkRRT3KN
CBMpWWZxKw9oQ6uUWcoHpWSsCap9epuZCLfqfbb6QoglZYeTbk6USaFMBrInzSzTA/OBjOma09Hf
GDQUi1yu1n6kzBuBhZ1zmhnOxmiYdG6UinQ1KOMo+f54UCaXgjK1s3b9ZVGln13GTzTBi5NcVWGv
D0pUDy3XDrZWF6112nJo8OQuRSv6weo//0AONbBj2Il59vG1Kr2SUIU2fUUXIzHGip0Qzjq43XZy
CMGeMijvo0Foe6e2zO38zxpvg6PdJ8/m0n6r4ClaYvsKFU/KdefGR8TfNqFuqEYFtH7r0uLtowJJ
h0VA7lcI08LhGqtvLLzWx6NNlgP3TAdLR0fR7o+foVQ0K6vLBqq258Bq7kFrtM81o9W2+9hP41GO
3Sn43t6KXqTOA9j0egCoVxf1At+th45gnh3N5swcbuozwOS4Isa83va33WmCDJxPx1dYtVbRRwh4
W0UMzRS2TPgUo1J6WbYAel95utfu97lC6d7S24wMDVe0jJJ3NJc+fsFK1aMKF0RcaVDvm8bz7JYH
0ec8MYdEH2nDXNLEp+2VbapC8Vt/sAzgkp/jW4X2zYW4+aQn/V0kKZf2+tqIIUHp/lT9meU4HuTz
w3jNPWNp2f1mSGCyUsHLE3lxgnyubK+beNbRCh7Q3yjtxuaalXzCeQ1bXzXQvR6oHQVeh+Xn0kZW
cPNCYs9M4syaTm1uOaAg551het1qBZDtA8rRlmedR83V1ecvwT33CxHhhmfzL7mf2uOGKeLUccof
emiyXvVWcZEpdyjqiyPtcB89FZZF2v2bNcX599TVlyLBcQssBRmME/U28YS90VsKWMtx/NK4hroF
qS/sY0Io1HTIbCYrsu7Zt2Ag6NgdMIV1Z5J5FvWQHPglLOCVeOZJdLktOr1UdrW0mbhQfiWHW/5I
OdA5czAVJsaQhAyxrHz05tAKoWKaQAToxOQDlbGq7f4NkVeV/Esqv91fGQ1AwyZq+NLFGhcidgXc
tZJDZflzt2mmbp/Y6RALM/AWcYkyG33z/S2QDKTE8QwOg4AkrGI9zuSbxS4Os/U0CTKCVDjYE276
qmcDC6LHERxWKWO2L+HmOw0h0U7WZSwxVqehbAEzwY91n7nS6kIcY8nGc22G/21czZX0zW1x0pkQ
iIcQwVi7odKj19pkxwd8FyahroxcG+zBkn2HQ10MmSb6iKw8O6oY9GBhJjtuPtiFSv9qV/tJHoaY
EwArhFDbO/oiuiv/X6r3avD24zVqizC/fPX5DamlpoPvGqppYKptlIkQ1WB8069QGl1FJcNe59rR
/12cpZlmdlG6/VCeqRsUCNnHtxF8KfRab81TWVc2qkCa9Ww+usfHYkcOl7dI5fBJuX4Yjb7rsfhP
XOqDPpQgzyUsRv+ve9hdWWzyuJLeMT2AAQfKIch2cZhZEYo+mdvXZAvGCbm2T8Z+vr4s5yWR6MRR
OPmB7LziaVDVwnB33hM0zJGWPgtwIZhENITzJa+EOpjOJ3Iu6WYNMhnRdGx9NbuNRYKuUSylssMX
5dUNehdK2F/HbiJnXQj+buYfNrkHZNZixj5Z9o3aXwoOtvboB3VMQ3yhPvzq8clB/0mQm+Pk1qm+
xYq9kTWzGCn/p8XECOXWbOYbkz9oAJFCJI1DxwjuRbMGGUT6A3Yfhz8wk0CeqXOUCYLqPXb2O4dV
ddKJ+FI4k77BX65W6KDhfnpZUQeKRn7IBNrgrlJuSi/Vdl1pb9vsUjoP1l9P9c0rwSYml+Tbw9Nq
2/Rn5TBC7uCOdtbaHWgALWlNxbpaC7Hy8I7cLHGznI6nWHwMErGy7DSQ/aFAehwfGuP5gBMeQNgo
WrhRGNBONLfYhR6hYL1TjUFxb7neVFH6WOgC/W/coi84StCAdeiH6TysyPev+0FrSX7iLZ+CQt2U
/hVNrfliCJoM648AaCdXXfGW2abN9TUYy9hXiQpxwzoCWYATGawd9gjHhm7PKXdkPgB1jnPXIH5+
nd6sDNVnMAnnMYwWnMnDIcS1+ZY0NGTkWTWb0N8d7/3AhUotNqH9XJJDDB53WhqNQNbzzOfMYAIq
urv2+3+HK2xBhXpk+1OWKoUMkH0YvLMJ+QHhKDGM8+V8GePQ6JVkTNyXu7E6z5rGJPdSLI8IPuX+
Un65qirwCqudAAWCNXLe90PyRWRLnvMGJtvmsvSMin7Ewg14cfSh3rNS1zNn2EBx9VslGXtFktq2
/CvycTOCukCx6cEkUerlMRCjDDrxljxyabiTQ24CLYJ9mMMzYoozAcHHB69GYkEePp6gXcccZJxF
4bboxxRwYA1Wtva9ChWHiPKma58hFcOjfWHl45T63N3G+3jETX/Dkr0Ln1k8k2+hzKX4zVkfGAgp
zDRbaW8tU1ZibzNDA1e74q/olZelI/G91VU8ptuBx1QUYDYnq74+McQq1NR2mcyknAUUkYtr0cR3
8cooUaHPWBWIyO1eygWXphkdSUiTMVP3ykBOKpz/YzHAX2uUVabStCbFH6h6HJ/7ul3KFAbhnRmV
JYLdwFAs/mlRNcNDml4rKulnfBMA6UhquXrK8tXkMrYKxadbaNHuUIq/cWtbwHaJqB6ymq1vNLGh
+bEn4FcnWJbu53WZh7yZbLQxpwXS+89iXB6XAbcvOIvCDUE/0aJCDFoNe2dSFVntyUh9xX4vfneV
edN2Sw53pfBnj5lMGVI/Z1YBsz1Sg4RKWMGplsxUbpviw+WCOAdOp97ru7U0q123Trc9BODa2SVY
z9hEi5CresqlKxImTi2OKDt3WbuLNs2evWnrls4DcFQyVkyK+G3Ga7WjXTDo4oNsdaK+HGeVbD1A
QqsqrFghWCSIuVuVlmSog/0lfK7W8qHT8Ps84J08i1cmdoFYCMJiLRwR4aN2Jub03Bajg2rzOE/o
ikw3wXF4AzNW3HyDzD7+Lkdh1OZRxIlO0vimua67EtTJVyKTJdeAyBGThXrDmCtI2rwkCd31UnST
8bBgQa0jGZ3bNBX/iWRghuY5hRRgKtfO+pwOoBKBbFPVPW6JhJ3xQd91bKWAHjrs2pYBji+8zCGG
SjTOv4I1CieBUv5T72u3mH4ubvPFJwE40JUS69HEliVVIdFmbHVpqG9qvOGVE7WnKjM44A02iaCW
zALYm4IgOGIVh4sRU1V184KlWztURZVt16TQYqPOgmhVbF2Jcwy/xpndp9H9qzwLKVLnlJ2bJuOu
q55wgrEmKBMSx06QOtVbihHkZ2BIHPzifTDcHVCjK2UYJkA+ArI/iTJ+9RcRshqa5gUSmMZRRK12
V2s8H9ZN+UK87ATpT/OOq231C8jPPXNZS7hxVhc2x/6AYgsvmtMfR+Ongy6nrw+WfKNCifVLro9l
LymR07FpdsrNqyt5iSORNKsqoo9LvSa3CsM3n+5dgAyqYJZ1SRXUvDwy5tyhep8UhCU0pcSgcFqh
/RGy+D5rD2U615qokRa3eXin0NnF6BqFBMhTMZSIca8d8jw2XLIljRBueDeLIB6kZEtBfIRaBKfB
FTIOEvW5Iuaa2VFAgBfpYlD3q0u1KRE4Xac8XmxtPepwltGyJ70RqjRLKtRHAmaPJAX5kb6jt0P/
uKsWEUouF+STaiQvxfAdXGYWwpEOUp1BO8qougM3f/qgTUfNilxccX0+VRWDeRAvZBgX90AjsYW5
1VrVJOcqvm57Z7GIB1AmAfOxuCIxOTjOnTKAOdBcU+zDel4NTpwrWEnSktlyMOu93++jGN561zWh
0Lepmi2SjjW9geZOcgvdXnNwzizupK8+3W28CZcbUPZ902U+agYUdONiWfcOkqx9aickxmyji087
f6l79HsoU6xARZuLdGh1MhbQd/eTFPLFG0yWabuEgl1evR+DvIhURsYtIp83KQ0P+0O3mKA8r+PC
PYd0ri0b2z10yFi66TOLSDa/FJuxc4pNmzQuFNx3ZRZQ3mVkMwvOm27Kphg4flqyGgvh3Ccs8Usy
+R6Tf1B/swlk24ZZpAFHqWV6Rq0elj/UxL4oFIkbODXnYwHdqJs+W6pRy/juLXFQEqptYMgT3XzQ
diMnyy3MjBt8khoSfuQMgOzYgjZ7LvoACmy2Qab73ZgLXUK13EBCDCH1jE2YRqmoB/9dkAZCZziM
VaJpsr0FGm5TlGYEnfDPmVJ/a/oHqnfnJFi1eULVPS7FwR0zsIbq55VvZO4V5m15LxynP2dTCTXj
KthuAl3h6IYCdIk3KjkCHmke2iCprfoMm9a5E8/Qt4vS9c0zZA+y6NbsA33oonj/ba2+HyydF8MX
+Z6N3Khy4rHnQhxSeswz/1l2Ln/RdchSakowFkGrSigkvkzOL71VXab58LKauswQKNYJIpTubNK9
pTP4rfW82DWR7aTmj1bcG/UFkVJI6tGxPtf19IZIy8hvzRiTSoo97i3X4hKMAS2PNjBSSt4GMSfG
lVJSLthQPyabGBZ3eFz2pW51g1/TLlygiS0er2QQ3Mq0XZLeg6ebUZn7S1/RqQqx/Ea3NYjikqsu
QABnkLiXmAtw8FQz71EI0Xr7r4qxZUn8OyEis4P9wOjEGuiTXCc7j5gNQUbeWy0ZqTNUXLzzV/z6
DuaNuzCIYevWCXywS45rMtn+ZjtpnKotBeSMzL8FLJWTNyFG3ka+ebRjEABh1s/K+dEvuDxEPPFy
ie4oOxc6AsRsPrGPXlrrkxjd0rSxmlhOWtawvUfEl1dNuaAKiwvg9zDLOkBYlFKow+vqar053OsD
CPzH54OVWAZnOpBxTnX7hdHMhvQ0RRaOFzQs3Qtkb+wRK8WGgOpaTz3ty8A31Bj0ARYlQWx2MJBR
OCXKdSfFsLxaUv/Z7nGFu/Gn7R6oyBVfTwTLvxc6YItF2vh2aJuRzuuS/nEOHC69xHAw0DZ1vYXk
QWJ60VC5xYj3zjox0TNrOE0GTFyLfvtgjH/rwWD/0XES3npwc0jfJP4uM5A31c8QmbI/eatm/wUj
1zc03Ll1iK4+erPQZ7CiOYl+kV1X4L5QrKNLIk85hOjrf5Gid22Zpl20YawSdZfpW/XjF+KSPqxe
5lu2UIP/B/VPzLnTcljDfAyZIQ+GeVK7rPsu3UH7tNffJTgQV6Ht6Pjxv4m6UEOYYiKVuLTyVRV6
uzkuqTcJZoPzYRsCunwWENFBxST0hp5BfwlaBYisgLlF5r61tExgTMbJESN/lm/jNgLceUDkBEnz
5ksGZ9IuegK8tCxyvtJa5zrCeig3xXnX2ym3FmSQ0fLiLIUUumCm8DX7GLSsYruz1jA4FsJ1dNW3
Z8iMl4aJyhIClqWfAsdMLyyD3bsEasE2rRmcg34GbsYMiKJnbTi3yqJK2vs/POapvXB8pfGomK+u
uYXrctNNl88eXiLhDk5WpIjpZ3dF78yLYUEAjwDbh5srYZfjpLao048jRvcnYtw/CHUbFs16ea0E
lsbF7sb5+LQgPqIj3XAIb71+BiT57mvFW4VM3lgr5/WDOwt/MzV71MAiuIqZgVmzLjKTc35TojH/
YtT3/KMjBnKFv3eBY+A4kC33wdW0kddHJ+4ZgkrrnSlJqFYLOwOz1pvkuUmd1Iic42SAEShcX4Y4
So4IDxD+e1tp5gP7b0rEFk8W9RxuRgY8rLTjFnxOTDJlEuoocQAbYjWNdW7Xq7bbae1NUGnETclM
XlNByCkNTKRXOLUQ8DChRCo0FPJ+/h1OqR1hFSwDJGnPSmEthP0geNKZ7IVYjsyBC1/jCnwLmTB5
haVeeX+MKsH1DMfXDWzDJ0vd6v5/clmHmqQLINmE0eZioUdEG1Lg9C24m4gxC3Vt0UEl/LaGw7MQ
lL1K1KGV6zo/LYieVgWF/R9xLqmlIfxdSmHUlGBTEjA54W/jbx14VDJB/Ji+gwrCAy8kA2vv9e9x
AMvK9RkvFvW7/hx9FLEp8Xpl4W3a1YBJTSx3ABIeFU6PeHkkUiTuX3eH7Gm9kkjJ39fIR0VLmChc
fVbw6RkkaNULLT5TYfLM78jxM6C1LVwphtI9ck5XAn6EKDP2v7UDc+sO2OLlukL0dO0a7lYnTB/r
ogB7edRtmabiD19xgDDm4pjywv4W+rKt+JcZWciVU3WriGUzZnrenxxNSHIdgvtVxjv9ImlNrsbu
UPOUMJ2lW+QMYCDxTocKKT8vb9I9O9wu5DZ5L7yOaCmKFtKm0kE2fXu6X1LN3mfbHy3qWF10f0hH
AFxRGVV2AtkUdAEWGpS3UJPhhsVcxsEWT5p2CLTSL/xo+VDYOO5LvhJLi0QjJ6tQKhX/7cE3LAdf
g0nqgprimnkbO+85fbJc/qcD+UMwDxs1O8gWSyeRHLoY01Y/jLTgt4KK48mg/3cQ0nEuZXwj8yRa
VvZfTtxEstaVFYkw2ZsOmYJ7DpVe6rruWvbH6xN2fcG8dGlFqs22s2P0lz1BNWdzuk9McOw6HJ0z
RTAIMFAmLmvIvZMdYgize+AUVNO6FCDHezVu6cnh2ZUKQXI6W6Bmxmxqf1hl1eTrO84N/NsvE8uo
WZg1cKrPtTsihf/heV3LTVBxqrKcDr2H/iMkIb3Fcxmhbb/HiqgcdnM8jjp8hNS2sGZ6w3bVzwcR
Nnzs1fDKhXqUqrag4ypigTbVpp/X0Eou/4RixBxvIeiluhQYCwkk49d50gQkBZhhna37mKgDW4tE
oHStILozgiu8UvHwQrPLiUVrr5fKbhrb6dgW48RKtilMa+2tOlJTrn4GU829I/tj9ezD1Md4y1+X
X9SNFoKghTzTPBMOgRZ5XRFBcaFZmfwWP6Ifq3ic1S+VMdclsfJOpMrz7vhNb6hn1H52zmu72gqj
s6ASns378dfdx54OVnTwmIn46W3xWBXm5hvH9qLMvVQrrGLNIFmcn39vroqVjBwfw1ubJljWNCrm
sCVHJvlSjVNCGGfazG6DMk7IBg5Oqjo3QIA9RX3EMdoxrJvsagFhrR/wX0dWzUtjMihPRWOdQ9zm
R7lwS+LSdmehMcncY2KRUeYoHLZIRoGQV+o1M3DdgHXkilpQO1GOxZz4RozOBeZyIs1bfl8TesQg
MVQwgE2q0zgCrNgsrY1mL9VZe9YyrBFQ8LC4Q9Aje323BxuuXBvfL+J21uXf/5fXVph5iHM7rct0
/MmYAeYrJFab7qs764oSSfqpSkT51Pge+aE1hDz9DWMtlVaWzwkd3BNhHvMzWy8G263Bi59kaMOG
l6t/hvFaT4t8pUnLVxIO2RxgZxFjfiukEjcLCzeV4L17aMJ30zAXRuFQSriV71Xm8refuQqjwDnw
oa9dKmTB9jrg75wPSDe2gQXG14JPpR58lUqUWu6LJKuiOoOb73U1NnMNd2JySzURAlCJTs/GcmU7
kFkQM64dzRu7hiS5qtdRSucOaK96xwI/XJAXXdqnZOLUa3CZMeeSiC0GWK1bUwEQ10a8DKKQ3L1c
Cgo2WTb3AE1zJkeKyhi+uVLVvNkQATe5Jnskmg5lMxWGaP1fTN1GGTu9G2yE58QtaKuju7Jqa+WZ
jRobaPqSDo1VcW7H8ep98WZ6KPHiQB9uYjFsS01GJXYRYWI9NKguaXKJERYhCligtw6osD9ZxEKb
O4fo93G35UTgNRGAX+5orrkL1+R1iz5/HUFrB08DXmFdwCyqyzEhb1yaiFnWjYPd7JYM+TcT7ayu
+cFc2ENvbAbmYWz9YH0wrwDBNuY1QOXkBB6fUB0fkOvxPi2+Oktu6JcQdmuEVtIbBFtG3mHtTv7p
hOo+iflANPFtYs9YYrfCuhPXcL5TI74pCMDoIVEPWvcWqvFHwMjfZIkFOLU0v+Lk/WOhlQsv/Fve
rkay+uxh1HW8qp2CALOEPxv6PcFh1uvMYi6egJKU5zcLDdQ7Py2NoMrb0GBg9MCie0u9aaq8RSiy
J0Tj1F7hX+JwfNDpyznNF/YKvMeJUme44/UzEtBzg297GKAq4BP4+xvtElNBbn3xW2iJT/kCBzj4
U35FVw6xuABH1RhmEU4v3vAhZwbvZbT8Qe1dOp8RCL8fQ06SpBEi4lOnJz8d+k7x31dlqTAFzjQf
iICqGc4VcpvNCciNXP4unpnXWGlL2awPpRglKWriSidJAGutinRlmcC+HbaokxQTXwvgJk8/gZXL
DRwDDH7nHVo/u0lDBfp8arhKI3ddKClJRCOev6tD8+3btAlmbPqtvXTKndtIa5G+AAPd+lSnvPbP
Ffwf2dH/5tSRGjBZWzM0hog+lGyyYk9TE/yXTgfwRdjgp+8hWEhC4T6H4sf8pf2/kvkMnukfcFsp
JNWhIsDMhJ/tn9jT4tJguWfXqbHoYrExGyytM6505Wl+FnDark54HoAfq6l6US1AsS/SblCtCiVI
3gRuY1Z8yj4AUJzGrVRppDiY59T4p0rxU6QR42wLjg3HzLyxS7pbyocDdoyt6Jy+gbCaO0k4Imxa
yxonisWKfKTaIxSZFQ3LykTAFI1EPhb5JHZcjdmIbwseuRVw5ACkP2UnZRM6EkncFdI5inHCypJn
T1aZltYJ08oGwD/ic4Lo3hpWsLMRS9quXNhmsaA/RNeYo18FdROXbcNMoxD9/MVKns2I7Cs3vheN
V47JK1JUCB11pUMQVl4DuAY68LG0/CycMc4/JxW6eYa5WdS8PlNMXsWq/AEieHhZel4SXz1Wdeaa
+ROeB6iDQkEtmc8fj2skmR+Blryt/jZ84caGLiiqyn371bA6wwp9YCnT4CDl9mYYeU1exhKM9FYP
zKFxULSIExdEB21nD0lsXgADBFXNZl7YrPFz2y7vAcFM16tX9kvgsCYdABPjKTMNhQDesuZjgKhO
kMN6noSCqnJbJfrHRzZ9huR22Pg88AyTvceDiVGh0DWwq+ysqe15ONP4s+lnIKa4Yu56WgSuI5gr
63sTn7XYMu1EW6Ce4qWVmHQB/uT/yzgNWFpnk8PZ2rCjD2b5Y9agICcfn/PGWfrskvxrO1ENBZ0/
BltgHJIXCBcikw8XpeyGmwXRJ8t1T6NcDoQ6FguWHHdcV7jH7YWdFbqcd4bd3yrEkwHBINjIi2eG
QHCvBn1oIibIyQu3OKUJ1ovsTtS3zSjbrWF27XF5z6oj1JQT+w6fvmD8yC0vRjrCuTmupBXfdp9w
oK+/+ph1CmUYEYOkeMCaeYLT2OIxipsLv5D3kcEZn0lpSSZEspjWASYaWwQWzK0WN7aJQ52AHGG/
h1RUseBzsRI3pssmHzWsuoUFRXlMRhy/KfZRmf8+OAiqCEohXzu6fRrlcGBIzPZjLppU1JvMeZ/F
Mvil6Vymqbnj2PndWYpjtl8k+eWpQ+q9R5+8fJqDlBrBJs79Iy7piA9cl0avWUToPpn/p0OQOXM3
b14wb1aGGu6DrdMjPgumU6b1+xxkHjjsu0pbiEcwbDW6kp99yG42NOIeeP6ciJsQXsHdJQaGvgic
z3JwvffqhefRN8Rc9CpH+eiFAFHe3XNgsbSoUw3x7M5wwgaXvVBXBe+fPCZgW/IDrd++nlY6q7Fd
vD8zMsHoz1lL23n695pbvohvagirFL44eE+gE6vSN/ZnBahaekfLxxG1cAAaSx56fvFEtdS2TJ/d
GDIZMw51MQx8lfp7K1imfdeLGTwQwAv4rArwLlIagMeqBVZlAHSaDN1m583DW8W18mxr1cvImrFq
WniHyPdC/XhWzpJKD9dP8qLANFOYo+cEtxsBi1no/nIAqWudxqUPEk7b8KIUxQQpK41ASzOt59Za
AzIeT9iTbzpUjBcmACPpDCVs8pBp0mmul5PK9nZEWuD9dLV89qAEiy+V0QD1oJNfp8VsiDRDys7p
jYoMd0Ai8ltQlnyEJQElFgYp1w8yrfr6tKi38vkP2tXU72g0RTR8wZSP8/CIOj6X2ny54bJ7KBSQ
neVlT4qOf5+1/qz8fGAUYYRqxwE2rW1G2qJP4WBht0bOVvYZZ3gosX227/Nk4imeOjqzc2mBmsTp
44DJ0d9WNFF7k/yWcoYqKF+JrT2OJf3gX6jg2c3c1MfqsP2lhXbXVjeQqMfPgGwjOutMWZK7HspQ
4X35DBqpqQLkTkIoKhq0BgRcx/guIgpRrkjkAtyJci7nNJVfXyWzOQwbLNNCbh8GqeL53hc6GfUG
vLJiEUC26LTbmAL9dKDqJGGCAz0R5Z94uQ6Zu+O25UKUl+c5E2UdPkP6+Z8xMtaqvQvH7McN0Ajh
e/oAqB6SRZThrNkQPkgdXilPSnLb324mA4X9Qarrt7LHtdTpy2Ap3lDjMilsDmEcg2YXi8z5kXHq
EZZPgmaj2uGawt7p58CM88UK32Bmyeob+K7Zs1VKozUjPFdgAhRRWPq3WGP0hSzMWbgs8qPACaWe
C2e3mKnFnmbtXAjOzoSG5TRQ91YAtQFy6LOHho9BmYIbD4YXU/BmWfpcGL/VkI6tYhqV3t3EedQc
n2Rs5EvBs04jfqKBH2WOcnl75RYmuHVoX3de6KJrBH+Lyay+nZ78wSPpy2lZCk78LMamBbz7nwPj
fOic9b0h9h2u/DV7jY7zdtlh3ksCX+fS7Jmi8BINgJ5EQlPedt7zqhDwfewCsjWaM6TPv42d93Va
oKjwDl3t8CyAb3lD4yJ1GKJjTHOehRADpIdR0DLtmTPUJiHybtB9HFnc7J/zZcJRTpCmNKUCdk+w
BPn1ygXo4+U4y/ak0OxSifP79X0gI/d6dOauQXCiQg1xpdGuMhnOwUD1YrRqB3jJaIY/T9jDCppL
xLqhdaBvzazpAq2RHtKVqtrCmFgcWuwLSq8xf2wCjWnzMtRBvjlvLkeCgdUkLDYQIswcwgkIT4Mr
ISqFKrG9gQWwfjVm3Vdw66yLn9A7seKADlZsC/isLRKsZmMC7Z78U+4EIKOyZNis6cnHyQmfnMtU
mmTGbZXQm8MbIIOA971h4f2G7jhPUkyT9hO6v+ePcJcgSHbQb9UHKvU2N17s/kN1Z/3//+9STYYm
7RlSI/dFBDFu8R6UxpsXa9VeJV/8DnnmNcWGVaG0uffHljboOF04pUjDz69jbQZkWSC2yAJlm1Lj
2mo9qzmuWXkdVizUs0mGbkCchXWCVsT/DtUHWimCCLgdo+uTeQgR9EvyJkZVz1iy0SpXITKWdCld
vRlVmORznSomD/zeph6jvP23Ka2ChIAuYK8Yuk/q7o5KXjurYEn+fOXFTOd1TBaXvM8uf3ehCZ99
Y035qeU3hS9EebpReTy+/BZbRA1xKC9wUP2j7C8FrjVGRyz295Q6WStmiU33BPGR8udgHBwuS7Qa
uLmDfC8DGH7MaMXx+PqpVqYZjEYe49zjjCQ4Qukqz2pQAGWnaO4L1PzeKUZnMsyRYNsvhNXlvCig
eO60fT/1TFWk/Ryuc9LN00XcyS+NqWtXNqO34f0FPG7BNqiczJYJF0N1Dokl869NN8jTLCoRW+fd
r0z8m1Sc7dHWzSnFNhMOc0BytL1AvrWbc5fLIYj3Y2kSXNg5lrNOKBGJ/qbXvagOaJte4kPdpIX5
VrhOuH9Ylp4dB2Zty39/pCPwNUlBL/XE2Kdqim7g/URL+miengJZyh8XmUc1UcJ0mnZSzG2NcUbn
cXVQ2QjXNVCaiiasj9/WMxfw73S1roM99tTbe3xBKu3FYHg+yHYSqER6Ap6rCGgwqMvW8cBefwwn
NU3+nMsAFD8tJY2On3VpTXFR1sqROCEQilMu817OAdVsU/3jCtE+AmxBcpySb8YuIpR02+Ma/ObU
amR0x3ia6bEKySzvxhSuPNZdPDJGbzyBn+Xv3ar/NVzmRNZ1BmTtQfH1p7SMTmnuhPemKZeAg4/z
A1nNiXE+tFz7qmJO0CSO3Ia4DHdIETWwRjBjmYhD9dZh1lKXTwI5Z/qTLfQOjK0C2Wv2AI1whZMV
vARMhctXf1Efwh1Kfejt+R8onaUhpJX5xUa8CDSOkODIJoIrbYngp8tKjB1qkEkainiEFNbeSNa1
iSOJzMSB+7QUOVFkGAZXXgbImKAwdxabQBVIH1B5T9Cjfj2bxArzyiRJ7LZJMEsg5EPCQLEMiWTA
fbogIb9y6371buyU+OgxPK4gZKoElQhw+GPFyxNKRnCKQ8ag1lGi9VjMSCDQQYlHBWS0tfJpX2AV
JEPO0Q/PFnplN4oTkIETzUrpcOMyx4dzCA4Y2XD5BvA74I9voKMqOGg66Hj44TlbDtUjuS1ai//R
Qh+THhAg3igT4KfV9gxeBpdfT66zBasXi9gGg+AahQEbIYntoChNp2LkCMmNkvQbfpqmSU99et+e
tlZMJnY0PFmBZL30rburlqAPaMo6qwiqVrN1iGjglOS6u/JuSLXy/PcnVz/X0n9yEmm0qfUGgi1n
h7W0FyKow0zorU0MGSjkEv5DOIDFgDycHkVdMFf5Ol0VEboJOLTGuPjCLZsCfqvWY//SSoKmrkSg
sgvtPflyWS/3Y+7HP/JGqcRYJO0ZNcW80c8Gk0dJ4j9HaALANLzRjCllAGk80OCTy41vrlpM02HG
nsF6k9mzn9ZCsBPfmba8NRZpzGz+JRGtd1jg9p+tTR6LX17PkHXEOt41oDyb6afmsWtShiIUcOu6
34Q7xwQM6J01I1fQMSaZJYuRA12qCNA3JHYxOIAxP+KsrQH8HdIeln6lOg5C9fS+hQa4AJk7Azam
gizHlbw0N58bd8nV3NlG/fD1M6oM7SArmmvsh63qYydCYP8jyIhq6Dx84oAd35fxBPNVbXwLbnoL
eIRXEOqOnxL96fLMx1rY1ebS2kdkNUelOS1mDzkCgmr1dqgAGxlaWmPJZSMnOO+gektHWF9nynzd
y2mUyBLSgJbIZRQ8X3XC6NuyKa1yS7w7TYRn11lmX11ZQvXmRGA3yCeKA54uwuEf6cHWZAqDuvkF
zqewRYYRDvnjIGQ8qURXvddrvQeRWmZJAoiRgs4dzHbxQlia4L6j5wh+6NVuRseCJChOMdT7MTAA
ON9k9czZa/0LYP7HAvVRhmre+cpnLChAuvAwCfDUmthhA/XsHl5f8T0vO3ECq3tTgwvr2Mj4AOsW
Vs93jwZnyinJIYXizDRDaneEBaUyeCg14uRnUCyYTiozrzQDfDKx8mfdA+17ZejnKm4XRm047j9z
D8RSq9/9SERcU/mgImhP5AuBov4FyPUDWswHTBg1nFYf54uJ1xzrq469c0U9cSvIRFrsSuqiHPzz
Y3je5lH+Fjf1k7YBZY7qZrR6iXGLdU6UZDr8VZJTo22bzXMd47HNhOa51lTJP+ztFVdOVjP8fWoi
HWnWd6fhNsIviyb00Cilag8g95rbjhk8BARUKwAq9LIxDyAWVn1sv9KDCiGdAxVy6jBRxBWOE/b9
eWacV6f5y6hoA/4cVtrkkvrKqp9AGCZcizdKaGDSnP9PoUQVdhcK6HlrK9ezZ+Khs+F8uxDd9YkV
w7CpzHI4Q8vlmLXSQLT0rIekk6WqeFhJXzJePRfUhpdANJL+mnwFj6iHPgRRpG5saWp5jZyTL57g
4yNrNLV7B5DDb1/eCN4o23TKfwVGGGOVlp8xvZb7YPicEfPdV+X3aYf7yKBEAW/eRtBpT78MUtDk
F3vZZdZZsb8Jm4+PgkmNKjIsldAL09+9aDislcgwX7g1uMYFrv39AbNIrbZS5tl+/nwJA3D3GLep
eBjx1jWjBvNUomjdq++0Jk/Tif3PweeD6z16nUgI7jjZV3DKToruZ0u4cRY5lRUziKLje3uA2fWz
5KzmxGyLImTE9DaTBkWHV5RGbMPrZICCvHXJ5LDCD56gW1nLt2h5PotWlXTGC5v7dCsVYTISaKtF
Q0HLBX82mp8V1z4PZwOTwVJCciWh09Hzgj5OHDMc04JK7a4uFMAABiO1Oz5fCRPZbW4BdZguk0el
fD63NkjFujQh9QypZRYxALnnn5cN/W+nyJoUIxORZuNOSoNs2rkIp0qA5QiV+69TXOPx8OniEDo9
NDjFhzJ26xf23esTcXgAYWh12JZhNscKXd3pCKx7u8ME58Yg/2m3Kf+uFIMFds/q1Prq0FIJUyZ4
2EEMGIMhInmvjnVOpywUH6+xa54wQBbFrhHJbbdnzxyWzlRQCVMNPy6wH00xtuWVC0ZiTtBPFQ2t
3Xw8uqdk9O+1kTZaMXChUlLx4LoGjSfw36ykL4FMtGM5PCYqDJ69ZU4sq8glQec6u2UTd0RSlM5e
C1yY0iePHm3uGCSEm5vFqe5b3Co4Gpc3v8j/vIgDE7gXREBsyBjXi5NtLpE1YlxqHHMITL3VGl/z
d3QUQRze2PUwM6C0WYH7bEqdbvr3OGObTMwGhuaHRibRJomzoNvLlEW234BEJNOkboNj5RfZDkTa
rY5X5oiY+C2GFxfOlUOX5nxdiGAICACQ/9IAdTDORKAhjuMArus6BSTVkzSt5JwJJHCRl+V0Db06
vvPM717z08cXIkNifO9b8M2ipCEoaPkUMZ6Y96U4JvUBUIazCjO+9xTRX2ORgLqeaf/F7ilIF/ts
UYMb4rV1u6qzw32mhzWPuSQ+xxEvsO0EAScpWt3XbhPC95Ykx9DgyYaQ9Xbi/+zG6x2VLdOL+0Ul
WAcsmotm+FGCyUcgtuyCiktn/HKtYML1eoh6Yi3Wi+ncepA1YlvmVSh/Lw12gzo24dbtdiGg5rQe
aDamzuXfxIoafXpfCX6yGMjns/sXg3BNmyJWIwpy0RSLb3KDSB7G/ll5ZYGvqhN+moKjkXz9Kdwl
rYFW5Lu7pz/4P0xe3qG3Qa4UR0uEuMZuBZbnaGmf8PZyIO5eWZszxF63T2OQZGVSHie7xYn6pin0
VWel0wHB2lyuCDNSAbIu+LVoV9GV4+w2c9AiSyTfNVye36Qk6iZUCbSLYT/nCCmurapJIZMIcoTT
OaKzPCYA4xt+vj+VAWlXLLNFYt8EUwAD+/2BqZbDBtGb0Xs3R3fkzlcpWFb0Rdxb45Pw9w+efiLZ
MJ1nUedX9UYKN+UrGu72VQnRI/bzDstN2k59UuESoD8mVT+s9PfHQfWMptSDFGhynY/H8UC9+TcR
sQncHSOGMFVI3uea12TzZ1c3LdgsZOX8NVkoIO/Xq6tceIH2mFZQAlGzHgEwWuZn1d7uXbmnkhR4
tuftkpNe/zhuZEa3GASnnZ1y1ef51jvp84N0SSUJDVsPJGAM2lBJcbl2GXXLsdABX2wuBldZhYJJ
aHh0WQaNBVJZA9S8hWZcDklyi2boAGQsIQ6NtVfdnrFqqA8Yu0wd0kijxjauMG+RDffV+DxIc+Uu
ladW+zs60E4XEZrkl/rlu1cAU5YxLtifb3cCaBRpH7X7iowUgiZNKQD5xuwo+ZN1UdxPR0nMQJiV
UsrhkhrpAcmYUEzv13GfHZQG9oE8IPB0OHSoslSLyrhgJrTfq5L11clsS+q08gZxVH7E4P/lZTWx
3TZabZiKJFZ5tTwwv7nzrDNsHbpW0sPtJbGoS4Y1Mx1fmWtU/IQXXJ4Op34YHbj0GXIpSTQleCmm
owiZHhT1tvceJMTf2XyzSHdzimnymrZdiOmfhj/ou65loKCtZSEXeeT+ncrtRbklnRwGj2m6Sx8e
+XyZsqCEeYGAbRWkYMjZHxx4iXaZAUGCEIsR3ZoiIxRt2LGaGgIRm7MbLJcyyPuD3/qbfi5aoE3Z
zL3eOACeQR9oUzmTVhY+KYguSDYW1Qh1O9kJua2LJKgCT/l4mE3AkHTJWsyNwkTnkott/pnm1qLd
Ti4iG7SkWefmrSjOa5+JRNZ/yAq+SC2fNb+yrDnWmmWsupzFPgaO0Q0y3Mom8KKDtt6MIyJRGpBm
WVSXBtoTMrtpZIU6Ee3dmq6g9ARI6ED5RQZpnjlBR4xwNIhs1Ig2kU2yQ9P6IBRL8nn0f2ZQ0ek5
FdCvSITVYrmFsxRGPNpNM9YuFeAGbHaYLbe8gJgDq/xaBtESlqJX7R+GQWZm4/jP5KV5hzi5SwHd
w8G/DNtclTKhFgl0vyQmIPXtNhjD+IyO8TpGl+ljNax0AGx+NXPFm3bkil0+DbSoU6d3/IE2BxAg
AqgPUPnaOwXOVUxT9iQpUfFVnrYGnf3VBEhJ7B5a4W9R8yd+jiTazFrti8m9eMZ/w0x6zj02+JIu
ysSzaGQmSnXhgGM9wRIgU+TkoGXS2QOk+UNW/03r+HQ7d0eZq8HKyQOl2Vu/FWIpM42ZgiQvZv7C
wGG32LBTkG0LdFTn0w8sPHU4iUBpP5ZlLo4vmV2vlcCxhjPV87WDd8ozdaUU9VzICefUbQ6DemuK
1G46NhJCEDbx6qY3aSvzTNCCnT88sv2t+FC0/l09R6Rpc3hjIc/Cv8Ztt9mPnn4Pe7u80DHkByR9
SJmvLAZ7VjBbkrsfSdDWutlX6cjVKMWbOVFxlzy7rnQ3MBG1B/9auzAI7vvgatLmw8LDSevDto0k
f3UbsItIUMg4jMhadX+mM5w30tY4n4RHhfJIiEmFObGgV8jroWNlyc/mgqw0eEytIXoYSCOyJifO
mB3xrtIkWUA9GQ+fRzNVE4GuEUwtLJJD0Z8NbDRobhOcQ0fJZdqg8BXl5GFtG7XQ3d0FZOuny5W8
glhFIrpkB/EIGPUekSnQ96m4pBqyIenOUhKcF3hK9fYW+fF/dJ3UdutzuMeaFUG8AGh58Ofbf4v2
r9obOtIUz4VW+V44Ety8fb+Ymh45aBhQzDsM+xKBW6KxaSkWRS61sK7nkSodFpLpFPyUw5DWfT91
8WEbuUDxauzmd2vHFzwJ6ii7EH7dhBUU7H9j3pYL0LjW06+HzpqRoyHIGuoZVWBUQx2shKFEPyf5
Myy7iaHABz0J7dFcWBgXWa11fyiz56FXjN7/4ON9Re35oHCy8duVQQn51nW5yybame3XYp3qHuql
LdpbAkDy6NXMogmlfo0mCeASIV+CLs9LwGr26cyaTuydDHUiqW6hUBmfZWsvF7BAyXXzpAwX2Rcz
rw1SQjZhMTidcijhPG9DS5jQ/Wf0R6z8c42O338Kef/Hw8SOyV0Akkl6HC9Qh5i+MUI+x4gShm4A
gjWlH8b9/vqHg3T+mTKXj2X7hAeCr1Cgv/ghIajJvikaCmkXB4AdfaOvPBy+KP00d62fUETVEsEA
RH8i1O2ZDFa54CQUKQ32SAMtdwV1Tv+azfDfEJJQomwDZYE3Ve7pns+bdTJZmhhflPgVeBSki58x
i13GK3rvAgBpUh2oMyWBl71Hs2tkRi6a22e0TyBOsXXC0RkqjEnGZ5NKOlDEzv5C0iK0Z9mMsjgL
Zo2+HfogZ9Sl9aoqBTnzJjmX8USJ8Va8+7kwKkBu0GhlJIF36bmk9b4GouSIzsBpCZC5DpLQRQf/
7PclBq6NAUySu4brprLKgg5EonVeKmQd/3HHE0dhb6os4T1Jxkh0k2ic9SK3wLYgCtQxLNq6STgu
N2V8aT9zjNPlRWtVKhqoO7KaHJ+T/eC3EL3Px9l+5e+Mxv0y0pLMhJEYX1xXHp9ANcZmVNfecmYz
RMNFRCOZUNFMJIoKcfQi785k2ZVZ4Rkynr3B7GuY1qGFml2Rp6xJZ62nExgsMmE79x88ykkn+mOc
ud87txXtO7+Eiy6KIrapSfiz2Z8mVKn/qiX5AHKW5gvOIeCzvbHkwE5FTuGwpd3vWOB4uOAcgrqv
8pJRqX7erOJix8EC4BgGpWSUZRdpE8DAA2kQJCl5+wYzPDlfam7ECMlRf78G/kcZcAguwwpSiLJp
IbHYLGjr4ugkEaTCqZWjcxIOBqXD2ZxqG/sHnSx37SIeOGOlIN0GCZ9o3fmCgahv/pBtyDVbyT5Q
AhcYMQYyw58Z18uzxkOKK5p+J9r8b0uRPPPx8pz40+j5ymrF2E+j8uZ/GQG0fTxdQFwNwbZ0L6r/
xpHDRejw04KzE/s/ocrvrxR8pf/bhmj/TXqXwzOn0bITYeajW5AYkxFz7pYP0VU/GsyA/w5zROKg
+bAMfj+3ZK/Ml0UiK/Drqbp5nuJTzT9YIoSRO7VLjeh/W0y26kipNjVHnBKVY70ip9YKgn9YsL3S
nTGHwPFOuWsqgp4o6KFuI8D+ZN6gkcVf3jA54mCSTRalxKPnLcDLFHWSfTxtdoSySzRcp3PCfGie
uraVjWj01HxAEWAOznuOIrEiVkkGsGCzeA6BMAsKnfmNoe4o1Nrkr+XKEYIGTb6YOdtR2B8tburt
Zvn98NsX7iXoRDnlFbHpUJsrJ2pALa2fEA9RPKAzUTUMecAgGd2N6RmKsr5gS/GQdWfimEHM6Wuo
rC+Qu/CWfnNM9zlRN5fdCQk5gPie1B6om72s/OVa1lR7JiXepi/yaGHKVK6eXMlM8i0DWxcI/Zds
nU/JEOEN/lUhmPXCXgubU/mikloxc0AQJAAUn96nX7xr/TOzRnW9wkIOrLsg8zLjJWklaKK3l6Rv
5v7NwW1R2Xmu8B+LPfhbIxw8q+GZuY4yvucbYIYNcpmorx93oCw65viTRoqXb0xwCUiKsACn/5yQ
zUv9LwBwR6jvJjU/O1G9ToyVK4xV+yNBniGIKhSdd0dQ5BMGqcke6ij9qbeAEsYvPmG4yZ44PFog
h/SYqq5cIjRfg/1fMNk69mTdr5SENw8nYnmhSgbK2Ni+pn7BNmUgCwgcKryCcho5F2ENC9DuPAmO
mwQv2/JOrZuqfaldUw/XPfDWzDYaie/CqIURs9hHm2dOxA2+G7A6uE14oRnJXfVktvvA9nyrbvPj
QG2I2Ml7CE9IE+z3CZiWF+hWykeH9xLAUq9RZWHKCJcwigDMv8Nbp6xZMZjF+qHIFVpbX48y3X4Q
MmoNVHkBdbYcdXF3LniWIsOR0Fw5QR+im+RitACF4DTxjXYxDyww5mYxV1LsjGgN+INNXK8hrhFX
Py87i1rNF1RjiL9y9K2QsNqIEqKqcDR+avd67z1V8nIZ4QHAd4H+lF08XghUA+Gp/XkFkCtRaQ/J
HIma6zo2KZEvKdyHmkRXQbQ7DvwVF2PYY9eUf3wqf0mhvj8Yxpyv6vvEYKu+tOHH4UJT2pSN4qkU
4ppnDya4Eqpr2FTsdW61cyCwlmiRdip9/Ri4LCzvpKR9NsSw6ppbbTUdlRIir+x4K8Rw9/gaOBdO
2dloyem2UJfeh5Q598368HbqPDqWRtGh3FboXvR0jfh1gMhyG1s5EqK9YzTpREm4XV+6IkD2X80n
368g6qKpSLvaT7B1JMu4f0vlD1y+CC/Hrz/gm940aGqUrwtu3gmCY0Hg68NWIDcIZ3yVBRFnMUcx
PZ6A2s0ZmnDYMZC68Sq0vNZsPScFQUlQr9sVgBVs62dWt9hcpPy+7DzoKiXXOIb/IxgXN6JA2wAV
3hNC+Hi8Jq0gxvEFJiIrn6ZGZhCgmotEsCr7L7x6Si7XHpSO49T/uSgP3zxx5gqAHMWl4eMJoL8J
hABKBrAGHK4mwAoV+bfihNS0p6SxJH1sdMH4byk5sYgI3SiE6yWIs9xuCwNwn7M/Y2WXd/Re4uir
AsygOZ4EdushMb966PKVf5hsvo2xWJjdvuhJmmKAuwILNBOkd6C3FSXhbmjgGY3bIKHaGEcQkMM2
+b5s6oCV2/dXqlcA+iSfsiBV07KpgrbQLTFbM8ZqXkH5GtoJo7+gGfTVCdl7B5atZHkVV6zQZQE5
sRPlBofUYW4Z9kU2Lgv1jpEVOYk7MUQV9zO2U66aN/dCacZfxfWGyzix88MngkVjUq8xb/D+tUH7
UIwMTB4oQxqkd/XGQH7abPmA1xhu8bitkk4SIGS5xMvEGUsl+AjSK9ra5HYQO6Z5lvGvpcYNSa6b
cjjMU6u0X2RNT87T9tb5OyfnJ3yuQafM5KFovom/kVJdzg7LeIfp4cIRgZUU+WTyepRcHX32KoMB
0///r6X5NRvN4c6zPF7MkY5bFyyaaURdJe987az9LYAVGb+r2XWCKARdfci5gpj+hKl+PVmgHV40
fktRUMitCoLDJnXTAfklvOD0l91ygPgCoTc7/zi8QszaPYqYLUTLlh2tA4I9xCSfZ2ypzIdWQnR+
QVuyrGo+7UeQMclvarqvBf+5Ci2Yoabrd+nJm/uZLMPy5xiJ1uEkjZDm1oszRnaI3BkbwdF+xQxM
3TQU/jq3uD/KbXVAdwpLB3FgWSBK8hPzfNk1PYKdsiFwZXDFv2qn5upDGsE/oljtiYe4sOvJnbxd
rsOEvsfj0FQis2K3qVXuPWuNIOPbDr5VY2p6Nz7Jf9Maa+UMUKgnHx/hj+wM+LNCCInsdP6m+8aE
w0SqhQ2i2wTB+MCbGko/zhorxXHDn+IMjPxPwhoRp58rN5r+9CLwPpSSP77ayUkOMtO3A1ATty9v
lMRjwuyLKWiJfyzTa8+Eln/1s1T5NqOsgdR5+5KiDv0YkGebSElwKr2cE34Jo4ULZOkHaUR7XOoi
GXfuw2/43ZBv7KWpP4dvGov0p6METFxBp0pykaZm1Puf2tey3WxKn3tzDVzRKXE5wxdz9nL25tXG
7fy/NBE1Ovc3VzG98lqveAhif7/ee5n4u4Z2CUcmDDJ7UvN3EzgCnPgK9Q9mcM7ZDi8e67pUoep8
0TcK+b/J+XMUHXBnpOgNJTQvsByL6ghS/H4wCCPbJpH0Dhh6IBDQeG7g3pNz28LcuoPsN676LgxY
xsf9MxYjuFIdfTNck8i8N9KcCbxBCPgWnEozDXPJPYO+BkhQLIVWYkdNW+fAPGEmzZOcAGiXLFSa
23lHUmVvMvbaE12E8BgxNexSlPyv13uyRP+Vx+9+gi/n0I7Ys6v/BQr1bQIj0twS9g5BJTMbB0fz
Pz9kOp1P1tiG1qgZyXQKD6ha7j3filmE2WAjCueiH6mzY3U8fQEbmah2tNxbwC3dF4kk4tqrjAzi
RiYqhvlHFL+6Zh6Swr9C/Rb3p6xm0e5IQUYlLN/kEBHw7dTQFTUPwcVwrklMG4z5awntBoOS7FVZ
Y4zGXbnJjfvckhUCbs51WDi/IOWpp71fcWOepO9ebrhvfa/4vFUqgE9wiKEveBTywm7B7IXZuuZi
lmMZbCSUV/LvKAxtN7x3oW83DWpNlDS74yvSQEH+2maiQFvpqF1RO0YP3TfQr59tZbrw7idCQyfJ
7oxYCoQPuffKfNms2i7abPfoSHjykV54gZuuXMvDoRCHGedT1O86qLh86zgzq0183N+Q/bvZTzia
bX6ZcVz6+YoSUTKYabOq+yOhrQPWGKVd9D+DS6lIqOUrbu9vp93UlIg0xmAWUh43aw8B/v+y7k+F
hSV2/VVEfF+ygcCo5Vq23ih+/PzAGuAGvPPz8S63+YFxkgGdlNpisCDUcguwxAQiQ3/Si2X34T+f
SAjY8LC1MHDqKPbLPN1xmcBYGcfrRbwXJCY+uRzMTb1fbAWo6y+yd+EMG8XMyT5PCfZF8A7JZXTg
FEyBdSzYsDI2glrCnUj2UG9LttFyXPaVGe9HCY2axhHXFZ8c4cVUVNoWHcCAuVgxK6qUepaNU/yk
pJtNtrif37zpinMAxysn0uL1K/Uz+KFCf/1uWzjKfu7ZRFyP4L6RHqb6c/j5YuOcr0G4iQC/XZGs
3rguQH/1DbcaHa3EO55XDtO71rKutIRkDNCNH4qQYYjnndzQC6jYSSBMwoJnRoGmmfc8tEyITjsS
A/9AcdF5Mw05YKRWkb+HddJl6UlT6OfKjUXBqIa1dU5KiqJtUd67/AJx5q3GT42b+SJMTXLbkxY6
afAAcdZc64HcUStgOU1AVFaaFdkpuGwK01LS2MvWkAM3dfINH9gFN40ifFYRumwNKTLMsu62Lkno
I5D6xVm74oiMBTuffl6E+J/df6EoxDtXo0eVbjIivC7LOvZMFonQEiFKm3+oFGBB7lTjs1kVU84u
Uqg/HrQojAPPvPv9xiMH7UNH75rxujOYL4hPoH3+eYaK+sv76b804GJXwBg6KouFiJgwk//wk+TV
9BbVZvtnLFr23/jdFQhNyIgBsPk9jYXQAWj0xdpf3jf0qq6EpQeaKfIbk0TN37Eo0e/H5/zvNHb1
mzEmjWp/Y2fUaEv1HwR+JDVEZHaNWOJlHMTNXiF7XR0OS15xmz2fyOmi0ypCIYbelsC7ndimN8fK
51zBhilttu04GV8aTP9Thv/a+PmEu6OxXPdgHFOP4vqV++fyKiYkVS0l4CIsPNbV64RBXGH0z+8N
t2pvFk6LCONQdnIq5CfHApZ120Wdd9H8IpcyhkWLrAfGDrpwOR/SHAgNrotIKxDQ9cDWeVKh9bCC
kcofurDwbAroXdy9SuygUTkfsDkSTrLj3c7/TAhoKrQqMT9GDT1rcfO+sAYsL8IEwn/aHPfe1a/U
duBQqXS1niPQx/N03FsyvcaYwAXRR6z6etb4hX7wcuPktMSYWJyWeyg40FxBInBhsvg/pu5CLmj0
dLv8sZ+ibFSHpNSKWQnIJ1RKi6l8ifaQt7ebat/F2ArhyEzuJ892njbtqy5sE6ugFevk6cjmvMsv
GICDmDgFvTEfVUdGk1bOUHBblDK3ePRC3r3/CEAzyHWwaqiuCc8qRCJhwC6Ry52E3qsDQAdfHuSq
oSOIwJRKfivCxHSw2d4njJxoQAGTRgD9neLudNCdC7pzkEyujF1oN8cfCwOghxV7rJElQBXodFG2
1ui8zwgtQLT6KwsbEHZev2ZI5GXrHg8e5i3DWPWLhi9Z6CdcfxVTdPnSGQziLe4BSsJOdgfUlkl3
h6vlFcpLWF6Y6rwOXB3rzaVomJUXSgq7/uXNI0TMJTDYHYYn3J0COjb/hJXg+Cukl9LNY8k2oNmi
LuxBCTZOD85d99lt/K/8uImRi3VdsVy80lRCZ5/tN2u+/gA+lH98TAZ/R+h1ZN0i+9BEnUNzDRe9
6Feixo+y/37MeKacS/ndSJYwRBO5keHabcfYHFONcSSD9ruQFjfWMvd5xF4F0+MFCcDHjbGTr01G
X7Us+kPJ8YvjViQQilCrWqxZuFns1Q04wc8cAJi1K1OhH3m7vXQjdHgBUNuOiYf129xXj1LoWuht
3Sm4li3lCvTQr1gwgGomjv4Kva1jI4nv/1iGJX3/7VYGDAnjmRxksd7ScDvIGsrNWleEkcdnwf6t
L9ZeZeNAUuZf75yRhOmWfhPsYk5+fb5JHVvnz/gDuQzB5w1M0UINIPXlyerQrshQJcuVBWe8ODLD
B0WYeS8r03O2l2GwQgMZSWVa/xjkup91uYj7gyF/gkkd8ZBlhIcJ9C2IIKR9WQ0N0vVgHYD1aOLm
TQMoYnzJYifIYdnWYT9CLfN2uaeyi9zzpvHfZZ73V21vp63aS7f5IGrxcfvheEUKQRM8dR/To1r1
CixIaTduPjyetnV+J4r5MhcD+dMfCgLbVUdMWoe9LY51DV8ZD/NHruhD6SUbm6hwpP7krYqbfrOa
RsLoRNBS4vsgYwuByo39oQW3aOVe57h2bfOKb6fxOO9fk2aTy38pVxo4/WftfbJPw/amIKT6CivL
gM/rx3l1cHPrBEE/sWTLIMGOwn59hotggQEnGaCyZcbw/7I8mB7zA/rlAFqAPUEYRwHUj49bal4i
Uogw9rzucIByGJpCkPtet3Cc05/INgMYsRyMeWIvNOnKUONk4xp5NCIF7XkTrtrj9iJnqg8nJGI5
Ddp72sKX6Vf7CIQFuRykQDnVM8AXZHGYWM/ylXbtuWB/hMRpG2R+iyyZOYFQ9ApJo9dgXIQBlzIY
/IvYGZMxa4c1QivuslSX6o2u61o/hFZigyzqdn3vbLCT6KU9ouKNWSN2asIUK5/kaGlyniPBcH/9
jQrYmML5ar+wGww6ANgavemLaayh6Zk3dbkiIHELW4IoBeDRM5Xsn40akWEPhFzCNeAXMoPlgnwh
Jh8WwZELfcqB9Z2oRgpiJ5wAkw7x8yZxpnZnAjd/x5N6zN3WsrZeLc3X9P0p8RwejZFODocQPkKb
syTsOo784KddL2gae7s7G4E8GBvr4aQDcWCMnsZSLFWu8DQMK34B2ndpAcIySj1TxwU9MLoTCzgp
PNv5QmQ5eMkkhD2QV90p4GADJCJ1FrZxq6jJ1fRI9nJC1OUiKsIY4Z+CHo6vMslxnj28dGJWs1VD
yqI4cTS9EvS5+mlvhLrWfS8uVE3q2YGVeRyxJtd5nYeVDIMeyicpT4g9uNFTEvUVVf15ZkqXz66h
fD4VXhfFdcV6ObLUODKNIOupsLEWPUzkWo1QpHKRtB8iFaHh0Jr3rrDYDvpMBb+kFifT3BoOZ/4a
noFRNEIG/oSnzbP4GCp8TItk6AXNWC9jC94POGQoY80fpltKnaVC8Si1CxGcl8tpLJW2TQSpXPlj
LyMngIHdb1JvvWnJk7rbXSRjkoGaIdU8YAfpZSePgt9xxHk/k8HyGkqC0hJZwJJ28KBUUPXkQ7VL
EEFJWJ5EliRTPQsQxP9MhOtQ29u4vkmQpnCklUZBesvUBW8i7K/cuow7rHmGIS7gJ50EzM3D0wiY
jzoxx/nV04d6YgaQ04c1w0pUKLTAhi73TQilFmyHV3JNePwywvKJ+2vjVjkg7aVY5T8zWmke4RGI
8c2l3hcGcoeamrkvmT9bj/ULclcDivMEBUUsvMrd2JcEW0/UfM7lXKcYNH7h706SlEb2g2Ueoql7
USNoSOsWTGwHOX8JC/I4IIyH69WB0p1AOTmONFQ3mrZ+KneIkcRl1B5uVybbwBNrRj30qB6p6uRv
jQA03gCs9Sop1wQbRx46KmT7KwumNMHxN/1e1QTEE4YkYYrpCv1gDP+lJ7FMozZh/xgbrvC17N+L
twAyE+GgVg2doa2efe0L+Futk2IS2VWFYvvm4UYt2v+753sUMNDIDfcwpzP9+CADRwlnLhRTcj5A
vsmaoayYIupsHVOJdbWO+h+xPLDiCyOX8b6KrW6B1Tb+Q+w2exkTGqkww9/p+Lh+8pVAcfXnmUJJ
8P8hiN96Ok4Ai1mGXkEM/DpHZlxFkgcNWXj9+ZokhT4ovzQ34sbXEzCz07Ng3tJlUaYhW0COoDmf
oQvZelF8+vfDnxnrnEhPXla8rHcDntOVkPoAf8KsVXc9NrVLoyRLB+u6aWKuVre/mgNoMpbnYyab
AD8MxU3G6KI5k63owmnM7RukqR3a2nbebTDaPRyeVtZ3PnC3wODKZaIOM/sz3iBk+hqIoeH02K72
1+2mSia8IBOqV6gVTc108Oz8XItitFsitXDWllMwoZY8k+tC7N+JdFvXqApfpTX+sM7BNK8NJ5Tn
gMHz/6OTXhKP3Idf54Rp1iRNJVZO7liOnUlAHWp7EyeNtE4xkxHV4ay0MxBlQdVXT/RiZq77KM+F
+4qGy5cBL4MXFnhrmt2f77WaCGWucHOSAjLjkqUev7eS1Yi8eYiqUbqtae5vXtnLKftWnadJ2Xh8
SrA2rgdM9R3AgqD3HfuLpWNI9cat4BtiqNGWSsDWjQ1tXt59IPEXv3aI0bwo0OcmOF+BLnrG07Qq
SyD0dOvfIZZoXupPgkv4JJWU4XgbERUn+eorzJwSsw7BvRGUxgYtCgVnbC3wosw49XasZ4nZctZF
EaVlBWa2TrDF5OW/INDGVE2lv21Mvkg0TG4GYGaPS1kDIRzwrFaPZa2gQKv9atn+AustbqBxmPjV
Ik6imqVEHLHeGAqwHREbGhaNx95gR1IHbysxfMSsaN7DaJInZ3JxJedua+2yVno2wSWRKcWaH68h
HYl/ghrIAh/P1so+JnGjORtC1wuGdAdzFu6Adhrk9wKbPkqPrmUKDi26FuvrYg140VStj3bhcKUN
uzPUI4muT03AFZ835pEoRuqYtW/p6jo9g6UNM2e6n96zoNOzLgCDGh44A/J3r0Z2b160SqPQNdnJ
sMUYfMvD6Qj4jXENgag85uBLaYmBjSJpl687iKcUsHh/7WIM1ek/7pDNS+vkOffjQeQY4BQRIbFx
wG9YT8MnpHAN6NO47Eg6Lyxit0k1F1RLqBE52e5PqOx4Juqj61Lj7l6sZ5KwyKN1ufdGp+cub4h+
jLQ2GYHOA1RPW8iL6bbtP57v630jDqKwQs9swYEDGcEnGLMgRqks0UvwMR2Mktdm2eBX+uwz8bQo
dQ+6p4X2JLQQjxooTz18NpaGcO9AajblSgFx4GRGqac31YHYUQ2n1vzqt6HaEvl6D8K90KACYm1v
GZZzrzywWljrpqr4CnJEUsJIx/RCtqx9mD7LuYapQY/XwChlBLdNazvEoB1qsXlZiylKvEPr9VWP
prIgQO8+2xATjOSUxJFPRlSTz4oc5+PpDYJGRqBrqie/uloyFEq/cnah6PKY9M1NRlOXccsM9nj+
iB77a8vt5SRXSN59PjzwlqrpC672ClalkNMxakJxMcZMiZYV1/Nlj46+NPMN0WFoca+yR7yZsAvj
zo7ZZLGgCeBsa+ICTO3J78oGnT7lYgBYqZUAWrCWwIIW4pnz0Tz2UKtt6Qmgyr6S+rwDdR6u5Sjs
YSfa+0pp5pK8m+A523flfQw9wlHWFRUi0LP5K7l4H97RyYUVvutkdB0yoHhS9g399JL8Pd2FuGXR
ShGOVVsuDqsu0w+x6PDAnDGixwSOVKNDB/E9tAPr9LrwWgngLuAPU17JuQkZb+bmssWYD1iWuPW8
MtbgfkTvS3iET1Mkw4NqJctS3VHCieux4vheJ+vhRqd3DsnsnGpgrmWPhvikOg/04JXTb5i0GvRD
rClc3/2NKDmbqzM5aKWLRl6qzJPYK5Ong2nQHRrTv+5rMv01blBiAg/X06T0aH6m6qXxAwaabnt/
GetGSglk+WkCKx7Op0MlFjyc9AHVkhmxlTdsVD1K4dx57XmuoXPhADZ28GFCDmY2DhMmPzjEdm1g
6ZMhnJik1Nw1qTQtmjSNl7/iLYWt8Tofludz3cJYKYDZNMDCYVuAqhHhPt13v3GlWVwNCL7AG+df
GxIZSPAie93ka9WGg/6UkuZJJ2UKph9smAQRRjXErmjS6trLotwfoeEwaH/+apWLFEPJKuR5N3m5
KXc//DZ9sTpVE+5gXtU8Gulf/kA6kf95wFeOsCfoEff6oZEDkqqo6hNTYRnsHSq51amaV6gpuXI/
BdSYwTvXW1RubhcZFk8Lp+Bs8oA2Y2Dom/qV0kZLUKuyOpJ60RvXDrrvPdtT4+8G8hydIQZESsDi
T9lAnTUEQKlWhLq5vvxa1dV0DcmcLP95RG9x/lqIhG63FSevhyxc0lr5AfpRDLHWk1iQgbWI7a1b
dV0PUhu7D8N8jn2xOnvyBGMGL9XjJkOM0aElfUdd9URtBpNDsunWp+Fe9JRGpWB303tie771X1pA
VyQV1IHO3HgMS9DVtQu+Z9ngh6ojXaKW7dQuO0KaeGlrjYGEdeo+LG8zQGjR+TqkL3p4N/z7QeDP
nSuVFTgADfDFjp1Mfbj3rczUcxs39OJS6nK+5Wpr9gdb1pW57/9r0ak7iUkTnn67iO7tpzTw7p0E
wq/m9PHC0iupP8SwqY8/wexGBNL2JwDTD5OHyR4SOFCzAeIp6jZT5EiAAQNYVq2NReE9yIVCx2ej
TURokJ+turc8f0rrUNmp4xqn9ku6rRkm0NPr34zJqeLAtjhfc/lNtsZtC64FA8Tpa36qrHz9gbGz
M1P5BwAUmHuAmr2o1D/i9/8M3CH1Xwg6dCb6KEIQ8eI+twJii9yrf7tRId/q5J+Er4UbGST85CiX
le+Yvo6xyoUI0fUZnWV883lNyuTYAxmQw9D1o9GoQrqBWo8t6FajAwh3Bzk8IPvZUwwxlgadGbq3
hRzF1Eru/MocXvVY/pjAKvYP3eJijjaJAr7VNSivFH+dJs8kXdSxmeWrxupZ4jOmbNeh7I1zQKdJ
/sAbtmgx8po2cXDWeyLCruPBQdJpL+pNZO51KQFFqWGEM/1R/iD2TNmqg8UTTvaIYG/rjZ7cy3py
IJD7UVgOy6wgQ+3TuSJtnBFQwro6ELJyyDoCPzV0TluHA6AZMRJhFuF5lX+ARGoB2o08SAzphncN
kSiTWXZRL2DJTgHHME6K3yJPy++dd/Ki27NIpBaR4HYOOoylcvGH6CwQT+2LLFyc7ve2PRdVDyjA
Asykgq1DpHObzZ9AkTijA9HBNyuCtVyBLMr++S1pxaVasWh+wkOPAaKtDT3oWk3LlRvZX7hcqkKs
NX3hojYdjXvYcpy0P05ltPsfcVqLm0KT+Z93xHc2iUEKX8+aIzshw7t27z9faPNtlrMb/d7I36MH
thjPbAs4tgsqiASBF9USglNN75B2lkHhI6MwYiT9kKx9lQHs5mOVuUZHw+BoZ75ac9iEd/P2hcyf
NEPb+Ut62xY3DXhE0GQeeEQSjnk3gjxQF1RMePKaOXKCLdu+9UxQ2Pgfw/WgQOQZWp5Q5uZCmNtK
5pGNfZVFuNr1vCXKUzRQnlFPi9Vwzlu7Hv44yO0jf34tFC/G1L7kSHuRZWYntVXDOKi1SZgIG+nM
97YjeySu2oT2F+1zIsxv4EZz04yqbpNt04aLRaWSVCXlzKiZc/p7lJyc59sjRHYsFs/2oOicZFET
wSbz6e9uj8+MvNaTeADJ1+HLFo8aQkUoFDC81sprvLjofyoU76YJWRX2hUFhQ2E2r4eilwXXT9Wr
yiXvXLPazbdlcqt9z1v9pKjhz49d0pUpnUOHdz5WoxNKW8LlNaeb/189hyNtqUbIEtXyzF0ZU+oD
CxJI9vMRWM7r9J+xBjhcefmfsj3eAJ+XYxWX1svgguD8TLCUV9uulkJqZjrhe3bpLLgozIFq5sF0
UFiRWvS4hT3tkQsYzKhRrx9yhoyCBfVi8Ys+LhVIVad+4o6gyxLWfKA/sAPvl39vHTO1h9Mcs6bd
rq+lopBIVi/OYqoru/U1Z0U2C8nDIgWu5rYNh93hZ47TOL0acjIeiApnuPNzbdpqVItXFnXifZDg
+f20yhKvxm04DpHal82WcHl8i1E82Xulp3hOn3GU0D8aC6RMP/+8srLhO2WMAE7pDvNkNs0sDFuh
mHoDJTFlrWvb+LKSg+c03S4Gl2C5zVFCIFT9rgYBjaeTa016CI5RtSOdDZyptPOy4MCJQJqccY6K
8M+DtGFeJp/3aZjbGMZgKndLQC3s0pDhwgSXwGf2WHY35UHS+SN0aFoNpBURYG2y3FKHb0sofldw
kraH8SbV7/GO38f9E7uD2wIUlH0uxGyyvAa+v0J/x6NZnSGB/b5w5rhqBe4mDhSSodqB5qvkUpXT
pcq0f5UPZlBdRpLpm9SJFf3ZJdaN4OStorprnYGPeuLv2gI2iB+msqark/tbROVpHr6ACSkHJ3ob
PbNnOpUcd5/BLmqdE5Qq/tKEHRvHOf+/1n595hgBnt0BPeaPsgqfmQ30CadykkxKyhOBNsA/9a41
Z8c2bsPDRYz+cVYq9GqDm6xNrEQvb91U823Pxmk+c7ZS/x39xpyG+7sakx969PzbiB81YN9NAQZV
jCTiNtfTXIdcTjZ3n1ou1TCHMpy5bQZC65ygyAb9vQhXotfSZlIsnggXFF9J3QnexInQhQJeRY7K
kGIUlvqLXFFd2ATM+iLD5C+tB4RIYIgY6zd1clJ5+z2VP502wn9wUsAMfa2zXbfAv6dS2TZjjiRg
WCt/W1e+ZsAzPXSO0YcbtOhbo8lVAap21lAeoirctRxD752OgGk4wZgh4/aw7FwWvo/xnHXAVj6N
8xwtmVFgfAmNoxc/sJAVZnnyTJ2w5xRZOwg3dJjBy3o4SrzyANiGETWpnvQ/PrQeBD4neAa5KiAW
WllTgzghu1BZIKXEUgiSSy28uwWj5Q3WQ0IBPQHlWGvPO/JnVSfSOcJlx0Ys2vGxMzET2QVciCvZ
AQ9n0PpyOZHvvRdG18VsuIurGnaEKeI3tUT3r3ghprAkFU5ofMTT/VeJC7F9Jtb2CWWXr81K2M56
H1eHIcEVMogYwgSLagwvMVdmo6Gni0/mfaASZLwFkhXNdeiF5Zg2GOs8yBPuiKcMhPZnnRF1GEzO
oKcf3EmrPt3nByF3CmFuGw0j8V+dnrz1hrZwcNHge87ohnU5VUaNGMdCvuapv0akbACDBgC2XNtI
s/QgDGQEEv6cU4bAmeNULB5Qdmpw+6VTuxHacmm/30H3wERa7mITkVMT9xXEHiJr15GXoN+rBc1m
UirzNAgV94iFO2RmYRyS+YQI8c5VrO3+fRK4Y47SU0fLsMde+3cTbef9a/UAW0VYVZ9334l6eY/I
xW3Y5Jzye/VMOzcgQSNJy+/9/ygatyu56zqJQ64kbTzYf+PY74Wsel6LZAZ26eh1Hg7cnfSiPVQC
NkT7CyBycapyY3UTlmmags3Y+VRVMuKRJDPb8un096SJt08FsIZw0jkdbdCRvim4fpFAjY8XIL1O
SRbILaOVuJ+o9fZ9u8pbYijSiFjR0l0QYeYqbcrid/qKoWu+Nuc2G0bVfbhBt+hXWUGCJg93YvYe
MmJ7lmXm2vKRLPebMoAN6rUrNoch8aPiV9rbAjxnEuhWQoeGE81nY/LSXvLNB/YaZGnWB18TmhRe
deA9K8anK8aYY5OjIuElicXW82rqOz74Oq73hlZZVAYGB45lng6E6nW22bJP4jlq4WHi8YuWplUG
1tBzA/I0UbNfv9772czSad/LcjdMYshbWocvQnM/blaHizNHZctMUhWLy6wepn6+o7v/pvfkF8ms
3Q1E8Q68LyNQh5+Zw/R9ZJqufgqPSgDFuDxy0rZ9eZZZ8IDvutZmQE1VNJ/TIkfZ2chtbl+cWotS
SLV6BP51pEiEv8asuqfn9yKIWLJrrGJ2605fifhmOTcxHjKiBwsB9tQjUatV67FGVErp/bLOEojD
6BOHRxVEDnO8PFgs4RDtHQgwjlIq4CjqQk5scobNiIeMmzPW+1BRp+FK+NM8ogIdJZHSOVcUbtEK
gjxKEI0pQjPsPst/LVZONT9bFvsGYPgBB+ZRvNg0IaaMwBNXBwGkOBebz23pfQrdF1IaXNVJufHN
cAfxkmfrztWzulhJ0nILJA0Vpj2baZGdCtoSpyo2PUw3m1IXL7qam7RLdOajmvUOGSv3KpDPBXin
/9YOvfaMwqyWG6+eEVcN+FPR+uKlIv/R4WfVyG2cxhji2VHuSfP4FqqBXlAPtRuQO74kZM4hdQVj
tDNGiO7sw4RX9wfZFfV96TxaxMh29ia6SRQiY3o/7oEbcNXtJFR7EZb33rxWNyw7zoI4sKmpKBZM
bsNnh7VK/e1oBwKgT4IJ3Dd7k0K1rUjKibIYoVZuDP92LI/TIlbhy/Kf3awSzhjLxiP/Deqcncv+
xFCfArTcOzQs+uHDoj9/40M08hf2NT/VXJunZiKdI7X1cjPQMTodtiasr9kgN3QkDuTqbGqHPlPQ
K8rT1Whtsby9q5o/QFk/qykFcnJvUzDvWc33LyPOzcdScK6dGqeruv4Zoovf+oW94oCCPL1QYoIX
WulYOu3ltT/saNtSKQoGPi4+5Y+jWMPTZ1pecRDlBHO5uJ34HhvDUh74FoVwYqaDeq7vo3TCq+hm
h5VeaK0nRWhpu8uP4V+DoE6q+hw/8EwrJflwHjRJupeIyMr/44WWyW+Zk9vTCyQctjn3XB9/p03g
HDNRmGERDWlgP39Zti/XH9IEjFNFslUTT0AIkHOWTlqJOmMZIT68PBmPh1VVL0N5SgU3XvHaSxmD
+2rk6e10sYNxOoOO2wNdFw4BmCYZLMM1AreljTF1SjazNyZ7u0wMGmiPA55Cze7aR4dj3DUZ+MBr
3giQadifDEQ9rxDS5ilEUiuei/+lY4F4Ma7Cu3awbgpnX/T1m0y8stDyJfhBmYbiyxCbG3efI4EW
LO7WUMGGzG3tbFa6no/XZRXASlMjXIq0dVGqEg1cJI+o2Xe9bS6KV8Z9/6wqYoVp2BhBmDfhC8Xb
J3FhSculkKkwST6aQMXDYZlHiPEtKV15s7oN4ktxByY2V6VN/3mFdY5w0LjMet1vhpDn1wAyvqGM
r8iB8r78Q824pXrjCF/g21tN18ZGbgPVPO6NKv9dL02eaZVYj+IYRpz6zOwY1UmsTBomd/hHqaEs
qw8F5MRb7z78zXkkcBcG4IXeW0vC2ZRnG+T7xVbmvpe4lZ83OYxQ2nOs+sBu+70mJZyOLYwBHLrF
7yJqJQdyhr41JjkgJxYawuiczm/j7tFJXyhENeyrlGd+P+mN3C+LHiwBwX6Cv/fwoEaCBb9RJY56
mrxNjEIvQuJ3iF++yzFXgDQ4z7V9QN1fwA+C5+9AgTCweLMohWo7uMGY/W/vtjKBKxPaIs4YZ5+6
emfFqaSMFF3rnUUm/xd1q60GHHJHvK9KFJD4lcxmbjmnnpFXJeWDDSQyOBZ5eb82aN6jlg0Hm8Ko
N6OnE8yYZ+Z3E2Hdlx38RRVUZWQT8VN9xNU+51hy99RvA06sL3eEafKgXtsdwTiqylKbVwHliv3E
EAG9QAquwCwGEnkOkTKHOe0AZ3RbWWq736RzjZgQef30/C+CF3zV+c/vDyoLiUm4fEW1aC1kjlBH
dLsUqTzwIJapm04ZCdCS9xeO7VlU+uZFplqMOpYj6thmPlVh8QdIsfpcR3gL22+LsB9RJLLuRgsw
ThVWrokRJO0CmmEzFmt0JZY/MH8v9iTXMDCMiuuFS9CSTdK6cRBt3lD7F2BnZ5NY+7ZJGYHh9jzZ
3LrZ9v6y7W+nToMnE+JoD7DCLZp2LjPnPqikb4GpCGLTk8G+MAUbpGvUo+IwUpEH/YkpAyrAbBah
SOijjFQNV4tKzY9KBXXWSJsyErTFHo1/toj1LFvFLrEVlrAfJbPw744sG5pmYPCOel6SR1JYbZkU
k/lFaJTgEfDoZ4l6dJ6uvCMFXxksIypvZoGGA18VNKxN280eWJCfL8ki89eqtHo9IKJHBIkjNKx7
4Eox+ImzcDLS/ZCIy8M9zLruT5f7Zpm7vMVO9nGKmGgtSD+m3ohnusFCOqaysj1LdqHZQ7Vyogw2
/vPq5eeIV1OIsI1Wo//Bc1kJMuTFAleHYYWwyxBvux6aBrtIuI4zuo92XwOTbnJE//AWyYP2cLoH
LbvMmaIrf28C/eF19CU7JxTVwckj1EiNVvFs5yxxPxwl7QEDHrLUDlCjfGnSGhI0d8rbhMXzjcKq
5mpWWWcN7fdXvqzwNhNM0CHGQhdymnE6uLO0EwpTuWnuRsRsH5fEIqP8hO2kxqHVtci062XS2I4r
EIM4hrRgXoZlpNgxPCLyA1BSZGgWYE85IRMWI0PQci8A2P1OuZGdfLUS5uOycKphwzkgjjo4lpOR
/c4HX2/x47B+/5DwhqY23z/WL1GvAuNGveKdIAI2AbnDlrmHOIFReu/W3mpuCFcUCGj+xHpbF2pG
dpy+jaPylPyumd9IWBu7MppxiK9uMqiyyjjap+oyjBmqgFydY5DKxQsuCE32FGsmqy54p7tKI642
Jf8milDbpVVz4cHaH/lUM4xV8do11IMq182BpgEgvfP2UmMD9ZczEjdSxuZWM1gKlfl11YgO1a+a
mNLdIdk5AcT8+7eG/bycFflhb14KyXCLVp+D0HUeJSEaIZiNq+4Pn37gWs4Jx/T4kDZLUfIuZZQ5
gPy/D5xy5eFKtxxjLIWjgCaZQ/1lmESLtW7gq98pFmx7zElSOkFclNRu9qeCgILiV9VceD0FZ2vW
EsjiY65dvxPYX2msztmedaWi2iwyU4T61rKgyq7dUlv428DNYDb0wXDDe1QOOItJdm0NFBfy5xSm
oJJxVXXJLZ/wD64G+N0l1pgSFqCMGSBz/x21fjPReUP+jLs/hPTZfrGpcaFRPqMW2Ufk7coy4C4y
JCT5rLIQT7E44mNglz+YheDYtgHPbaQiLtWP9hbNA0gmJV1pIdS+pZaaHnSkKpKIfV6fkOubUFLj
Y7u180Vdlj+rweLHVJrY0XV4B4mxDANbG6WH3EgSQPH30TmKUtrk1vFdc6HTObln+cSImfrB9jq7
nPAPGfXkk5xkMqwI4Xn7/R1JPBfXqZbR13KZXiO59XZiZKiVdxqy1QNIJ7MbvfU9C2Iw6DQkCgrY
uwOG1qhFOF7B0pFx6qvfZf64n6WDME8n8s8eDkallgTBhEeaAdDYlOG2xIPK/dpavsNXeeN5gvE5
Y6zK7hsrDJY5hzFrLywwOxgK09dZW6EZN6hYcT8A4pUNPMN5VtqmLBepEr0UdmqJCi77no+xyiSl
jrDq5Re8/wnJnys6gKlAeca/sv5qLRqb08R+pTzTzPuYSr2HKJu0AukStbSi868XpbcriTL9d+Xe
/GvfFc4+u5mbhmhvJQmKamigLigTW6EwR+TN0H1+FgSCRa2ooLxURf9yGN1DyPWZp/rdu0uF/Dc3
TWput/rIpdRwDk9m3RzkypvAIk/UhlJ8cJmQXe+XHsK6tHADNmLhhnV0CUxZE33EoX61JYgzCeDI
X0qk1F8+MamEYJ5qgZVY46TadcZ0peRoj6OkTIbXhRv5qdlNUskJK2AyrSA3sLjPwIcz5FyO1Qj4
Xy5kEK2xgiIpqZswxJsfe4wtfcXTtNy8xVumuSEndTQdmns1J4XpPKEWsYyKiHIHUCxp5KljSvLz
p18faPdK2TcYdmhKdeR5/hblmszNPiPgNNZoxgLkJj4742FlNeO+HJubxewwJWOa81XJ49qBTf7m
b0TpxjsygBW8hHjCF5aqsKLvs1MYq2bi63SnkBQK9SoRKQ7FIL5anPWPmc7Dvn4PcUOx0gDVHYnQ
s/gdgfvLT8ohRfbAtGfA5joXqyWo95Wra/7iNqKCu/ORiOPN2kwh8OwwJwORDcpSHvfQis+Sm4S+
lx7br2cX0N8cv5CMW2LXihRF32AqyRPRyX0gKN+s49BM5AmsXyTR2e/jbvrGnZuGQC52yslNSUTk
GaHX8HmLamX5Jn+WBU/Q4QV27z5FReC5xDck7mb5m4Vozj1y2nmdVJx7gjd0pnDTTmF3NvtM0UKv
ZRkS31MzGKAWrdH2vGLIcLm6hPcOfxoPIrmmG65WdQU4Ydz7AXKSzGxd4ME5EqnUrcSPUKJpR7/8
NoAGZicbxuluZMwBpJJLMNt0CiCGMg4UqUadxpkMmfghrwxXpjrRZq5lR4vi1KIrLIwjbC/4zB1G
Wmzr9prk0nX+3jx6ljOiL57LE9QjBMMStdL9d6zsrowJVtlhp5C1wY7PV7ZX6fzeAW8A9OoxdiYm
SiiejgfzfCv99dTg1+DosfvSWh4FHzar8zXEET615XNF+LfT7NQcthZ6NzUrdfO9fjbcdkbQlb4f
xV6JvMGZodesafXMBewVh+pf+lhodnirVqSnyp/m/4iqYLwJMZ9VuCpFvhzf2dp+LGhifT9+i3N4
7Wd9YTxj0AQse0L0LrUT7H2WC+WQbNuwKcWsuqG7ye4yg52PDaAlVpyUaWl5cu5pssn623gbLsfS
TrGZ0etkliKTVBdPsXugMGhK/ji+umXIlc4M/jtyKBSp13O6Je6lYBfL+p86IoKB/qAq5CrezxD9
G1BY7kGK61JvZfCuxddFw/wPgyNCNsI0sPkr2ha2lyrg+wonMhZPhpWTLCY9vBowAIX9f0Fl6YL9
q7LR8EwM/TXm0vHjHYNnPMU6QWjYDDfsUxYBSQggOToli7eMA/JQ1rlfsfd9yWAUaPV49BkKko/s
NJZyDHKLN0FoMeyC19bJUsELugwW1rQIFGjnxz3Pg+dZE3xe+3CWZONA+TovJ+AwoTwYjFenE29p
PUfJH17FvERr0sMDSHohsPDsZYXxC81yMvWYK2tFruEHnjRhc3axqlDn41BXfjHZH/tgn3bM4IE+
WoIXYEIgumJ4skW6A9IUqXsZL6GVEakrztlxh+zjk+YYCK7xRafuepZFkv3VNrTx0Mh883npF3PS
wZY2xn+EFaiOM3O3KH4xuOtXYvR7jxLzQ7KqQGrDGA3Nh7khj3xJqoEsCrPR2kTiNMUexTQFWaFg
+zXyd4+x4OOh28+oYKsTLWaDiMyuRoRm8A5MScBZnE8S58/kNFPmfICzCWUa+ctsAnW8CDlbCOGy
6M+EPLEJhpEsN0WbHYDlpJTpgeAUGqewlxHIBEIbtCcuOetp+Vxih2AMnTzQ5bMD8N+6lZP9b+LN
OcurHLmrAYDM0PZwQBdQkjtotWsNZNvmwJr54xSjEVIQNxSbQK+pu6TRQruCeDTTketI3du+LNZ0
jq0yIjSf8wr0XZIOSj9LL1Pjc+Eaw3mU5m6qXh/5Q29KZZahjEdPlS4d4B/kmOUqPk0BqGqg6qi6
u7IyWBdLUtySdQjBJAyNC5t91lJvEBSGdCtYH/EiZGEuWxc26GpP3Oi4Cf3YEA2DBURScjRyBHnr
QOubKRSCJJmQBMdZEQrWGHRNbDvFiAPZUNdBN//4MrmlHNzmag6Wl9X4j1dkTyi5fPVnkHL9QBFd
7V8laQ6MfeAvn93zqProhvd3JyjjuXnE+bjba4LUabjAVBFJT0uTPVw9iK10K9j/sKFfUqKhcWwO
xcLIWgoC+jJ7p9PgnI4zurr+Jpn9hJzDXBt9s/a4Xo7SxB+XkXqQklJqpdR+f7Pnmvhw6Rq5EK+N
N7A2RGLCbdmjkdjTrhr2shNe/zKaid/oULA7VaElrp+1jLGBb/4qE5WO1Y8Or4Z+K6dklOCLPO7V
Jw97vOxd3mf42QWZDPd2Vq6dtXHbBe0469LJWvh2qMinWBieeAJod66xUMiWTvkST7B+AvJGYowl
ZyIIej+mAwAwJvGUUspW6gPS8/L6ayz7VCK07H3urMNwFW0xtd6RCaHt+oVfxnsjEFjMDNHsnkV3
Av9xxktoxP/2yFuyQDTqPiJ3g/iJl7KkExNibkOMm9tqNzke8sSTeLOxOZIYbspyOyZoj56Tttwj
7qFmBtUwSSfhNnNYeGZhHADD1Iy7zsmVPkX9nl/jS/rEDcTHy+9uTxGEV9JEO2XdQe1uEysNhGyU
qymNDj/7zh8emAbO24NVV3HI9f/Vsk/9nB+xisQ914xfPrPHwSUg6WNEnTOnD4pJirgY0ESOWxbk
xOVdgolLLw3SVpcLjk3g3k0HD4FfJkpEEKJ8BZQNC1uIpXHjAEiXu0dw9vcE2BDqXgkyey0FfrD2
9DuQkmHwrSwY+eHUW9GujTcI4T69k8pbvXGOGhtbzkyL9V2zMGM50BoZaD+/6VdlA7cSdXQ1LqSu
6HksNSvAjckO7N56Vay64JHE/PLSTWL2reWVwxsO+POJAhxn19BWiipAqlpkJ5lhfhtD6d16x8lN
ZJpzXzi614u8I2HUw0mQ6c5hVySSNpIa8+vb+WvbudF4WSIIDVQNjdAtyngKNfY/a4dgMD7secz5
uVWOsLlA/gk947EUS0STuW/J5lDMAE/Pw/5cqnLxlMCfWKduNCzgcMm0W4tX3/ch68Ly+3vV4c5l
oY59BCqeInUJgAhxtG0nbUyCK+UXIx5F3CbqEiAvWqLjGedARSn7bEsWeYAHrMFZrCkNU8Wqpn7H
C7Dls5gsq08qg5gU9eyVFnSsMk7p3m/rUhJ5oHIoO/vzoWw6U5+xLVil6QsF/5QZkMbyCWNZHp/F
mrc1+DJln7dAjgA0KiR9NqCuUlmIMOvV4gY0Y6FtTqXyuEcDyJ4etNpcCbHGi9S1Z2ZtEAXI4gJm
vVy3pOjtrhAlJlwPiyUtRNlrr4TQvwwUD6ewtJiscipviOlbVBD/fRvszMyzrxvwMr/16GXg/y0Z
T8mqM5Jt5nC3sHZjcdiEMxCrGUvMOb4+jW/Nxiwjfy6O5GbyMahHahZFvQ0hPtr8h5+xV0TrKUeW
V/PfO9WKXNO/Hb+CJwQVBeihbILo1tTBbEdN3yJ/DwnMkvgNV5R8ugjkJu6rhISzdN1OJCd2RN9l
GqlzysYUstwHMI4lLNWIGZ+nlALjiW/BtvwF3GxbrH5xKqPmJAESKHQL9pygPPQnG66sTPiIGHOZ
7A5tOZd8DJw1VQ+YvTX5sSNwOtaJEgR+uunG8WI0H8kodbjTnGWjBJLuEuc3JMIdSAqthBT3TbO9
is3IxxnEXns7Kbil3MKSWMcd85ggBmRUxsDH9GNFpTRtGdgYXZOzNjf+FLm3SDO7/V5L+KJpxmtP
lPl3QuWT3URjYMnypDHVmSMDZG2EYAxhHkZKfjn2ehU1+13qIFOHY58WUf4x/AtNMy/xdPR3b1hR
GxJrwejTh2jRAmbJwsf6ehI1UoYXlwRCm1qBslxlhE8EXoPQPLVaR14UBzuLsPjRJKWV6uJJTjCu
q2Y+Qerg5M0wYPplJ5cDHp3UlZc76iUyJzbkYfFnBANWNvC4ra6H27Z6Wi9P6qn6iNOqXR1078+4
TxBXxyCDT3gtJs68jvE3bOUXlolC6TL/aDe9NnD1paDq/6u9pAO0RZzls9jS0L0nSc5Abycf9eby
KLK+EgAlYkYh0oPtay3BcwPLqcsHY467v6PuaqrWcVxnpaPsEJCZbhoF/oReEeDgf3ICwg1WR92h
VTh6nL6n1s+KgEeTwHaS46gDn66Kv21SqclrtwSYI15kIDNiKJtys6V3PnO3Q+eE4YL0PHYmlAKX
MuHp/y9bicSxBXEtDJHHgXtDm/jLy8dFrp/r2klDQr25t5h/Glm87koNZatcO2kS1jnyt2xObSo4
6oGrKJCMmxKnSgPiW5WO1O+mxPZnhqEMNFQFQNSd3ZUWBjteyNxBXMLaxGVDEYUrW0y4OV73efvY
OCD2MbOCx82UzNSA3iaMQqy1WayQXm8Mns35m/pipQJMsI9n1SvVyW09q1joaH1QsBi7tgx45r/W
Az+MolsaZbMqPvVj33VcBOFr+4lx9Ja5ghgl5PCK4/nL8yyh0z9MrJl4ISxZpEkVYkt6DFRK0kVe
OUfrjN7X+AbI14ZiW3QsfG5DpUAxnnCF2JG8bgWFUcleLycFXaVUHXRAntIeNVwmDn4T4/MxFpCg
nRuKbIiItfWvVH5gHzphpQZY/WPuRCGnkHs2npIgmenyWt4HEXyUvVzBl8CsNuvzXzEPfDrHF06C
QObmlcdMZacMbUpPtrKQT6xeBVRAAIA4/HgYbjWtheKrD7F0PnTix0Q7akYZnvNuh6yiPP3xN/g7
mtAKJ4YdpVPjeruhOUkIKQUm1vCYpOsDbWkfU8Hgs4vXANi0LRcnPr8xvZSUorYl/QxSq2QPNvSx
YzJODno82U9/+AK9rxyTH8aoL9NollZw5occcqHcCf35kITbrQ/VX0Tn4DMaHSXI54VWmJrUHpqs
NhQ5iTMJ/qkv9UotWpNez4WmpxIA8JBPUJ2JJDy+vZkg1PNrLpWUKAbIOCD+KW2qqZh/KxO1hRnA
A56Qv8uoO4rhrKLSkIWkJ+Fz12s1pUm7dukcOfaEtG053RYiZ0HL4WUsgLZvd62aaCfKrC2esgqe
Ft3NpVSaXfZ4Cx51pcIuZCUtwV/8IlKQ5tNo5o8ZtOiqb/Jv9vXaj9B/pMvf42B5uZBF1vUZhh63
zymEdI39a9ieaT+ok5H7LOBTuSapGncxnkAKBlnVsc/a7UaAcUxq+vGvwck80pb/RpS7R/3N/INY
mXSlsi7p3IVsZkOJ1w3mTq3zCwRMlBPTP/4vfdCBE1+XahvbpVILWW/z2L6DjnqXFm0fQWz84IOO
tHci8QZpWBMeyC0VvGOYqXCn1DwgF+AVSfn2MxSNz33mGlc7P7jSPlEZq6CTzHSle6uA6hY2IFk/
nDSTrgdw8UVRxnRz8nhGM0vViJRggWNezo7ef7a97D2aQfYpreYL0mdmdo0IGfNR25E1wIT2GtlT
14ozesyD6K3tCXVgNP8tzimeHYGP5FpOY989SKlhn53nrOsPpdAPXQEeH5g2eyxuVwBG72WGmqyv
xGGl6FtsW5TtlJYj6Vm4NjSFjk8i8t/PsR/OKrKR24g/sbZZp9HepfSdjCEN/FrKhH8ks2B0kF3z
ycVouUbCKopKmT4I5wfIq5vbb4Zix775Dht+x/+BMNTfp0eUGiFHX6CEGmBGdedd0a821WSDeGxv
pzHmT/ZPb4S1ke+S9FQGJETfhOwJA9JLqXkTCYlW8kgKPgIO9XblKNgmltziIyp3lJ35Ij3WOOXC
ff3CUV/UXFIwVR4tIJ2VnEceTJWO9v2CjtGGEe96AzRi06wUA9pwKhx15Nfrt4tNKHF0oU/QZ9dG
of5sYANabtpp5tHIFtKQoEfkg8UbZ1K4KAzFIRWytXzOfwHDnPt3STNxb9fwZ5lCYxjA6xomtFp+
ilfNJrZG9qUv08ZjNdvshSA0cn85FwZ0TBQR+dIAoDUSn+W8qAldhZnNmxgPVQdxJMv7Nz9n/lZK
QkRIt7lnvfWnUeuSGieBEM1pV4xCiBYTHvwtTCo0fsB11LywwWyJbfm+9S9zFdLIpb13+bg/PWJ1
o7fMsRuLCtvVXlhR46OBgikG4Z5BhaiF0wVrSrG8xUVBcMWcFBlMLFEKmTDfeuYmb0KM+/GXOdhz
gdePuzBG8otNWB3VgciroICf8q/jQqC5bWZzV9f1bFPCSnWT1raaqwMeno9+UB4CRDINExqBzfgv
ZsWpXgvRlgG13D65NH/F4DTjzzCoil1j/FH1zSkWiCR6p07X0jybn6Ts+vTQ6UwSZAq/xW/brAlz
00QttMy/QgoPV3iZNLT2IGRWZCpTJW/g06zOVUV3BEUKPzTG6xWFNyKKQVRjKqTczo0pMYNRloVn
gus3qEJp6vmbWMpBystbd+wA96x1cpC7WZg0x4cJ4w9fomaKmDvPeswoLzf+bCXzf4GskxRmUj/y
nT2CEdLir33b5I5vb0s8RfGg8YlSHGYGZNDojPPHgYZAbxelfxQjlMDrsMmOLG2JtLDIeYys3Wkd
28ez8gtiFiF/svLkxqS/e+X0mnztWb0gGwvZz3NjqdrT6mMYbuKQ606/YRPE6no3I7dbhxYpMTvd
PMQs4PidzP8mWcVYQ+m+XtPjFKDDGjStAQIGh69s9yXlFF3JSdyOOhdqiAagBU+We4hGOWDlxBp1
JlyZ3lrTUAcHqRDH2V5dld4KcoO1viWagF/Of4+1sg8RQhFiQaTv4SaIRc0xb1Jl9tZzFRk6Ubf5
Oy50n/DCYhkE65QixfJBSGiixhhMgSll8jSxpbXC+cjOU2kdBeG9KbZbl3xNwsVPmAAGmkTbVXWl
asIL+GoWxq6GB3GQj9eu8eWnjjcA8Uyzd0643aKht1KSDWUUgxop0o1ouHvsfosd7M8o3GQrWNkr
+Qixa6nek20xRQaV0Y5p0MElpx3abt+OYpfSp45Ao6sfZHjULSn6MPGnXk+7/LYdQGKhzLmr1NX1
pkySrCjNeufq5zMYETwSylCnDTi1hEheLv3jd0q3vv3oSwTxVf1OHhojTFmVqjkYFhohl/2ST7zN
E4VjqETJzP6Uamvc3Ko2bY2HvGU7vWCfhVJfaj98+LpU7XtFj1JZAtQQxG4rAb5DtkJhe1RY+Z8L
kwYnesjOH8homSqVYxlrgMydBA/lxiG6xWhvN/ejwOWdbcmQYNd/FXJ6sW1UtsqbXdeN2a6zv6+m
1BM2MjRtiASLwqphzyCki6zLZRO376GahqGh/aMPSlhVwl4nehZvb7JDIR02KJmL8C7KKGdJvs31
H0nySKOrN116pZ6kYr0koYtjugi/x3LElgIKS6RdUDN7a9FEVNUzkPWgfrtNMOk3RY9ABmALqDUZ
HRfdF/9K0ZAElg69Cv3RIPLq/Nbo1U/tzH6XI2zW2ggeWZ2iNuIeQsvGB1OeaZQicbpcpubMGILG
DgOMS7fkoJuu3/35VErSJ6OABmzdpjpJTsupGs/84vQw3KV1tHWnVzKv55R+xJHTbeqPc/Z5vtal
HCVXTIfraHLsqHZ7lf1Ahhkjg7nkJcTg6rN919ChOA0XYolsFZc7zuuJeZ/AMwTjOs1sfN1Yrtyt
15d3ka5oXpAdXsiK/+5olvFIG7y+ckdAhyRfFHIDZ8YCzNsQb+EYI971+CmnxopAdILtr8Cp6/HI
kMYVAq2rd3UObnj16d0e98gcPSK32VY+CM4x05BuXeQR5ZyTUmxrtSBa9ze1P2Zw40udORbfDrwg
ZiLWI/kqT/VbzCe7yQaauEShRKbqGktDf1s8U+B8uWPFC5Fgi1yCnXjghg6MrwxMAmEl4v4Vcad2
hnj7d6nc8+IENeWkEOd8tAFVsmvOFWBg73XqmQSol06V6z22MDQQavRM4Ap1lINw8nHNN3XHQLVJ
9kuV76SlRryU1YdkncrPRfUtHgVhSoGlSeYBjsiP7BxvpaEZeKVqbEtRzaaL8s6Per69mEiT5azu
6RUiU8le7IaKi/2hCeuhRKLRuEGrfKPT6DZKEum5H9B0lLERl9laYXriME3RPuSfBh1OtkjEH9GY
hBytd5shYg05ozOhwtxwb97ZTpJtlFdier7en87zkolJj4KxoONWoT7R5JqwounWAmfIkKBOg0v0
CcghTs88XH2yPQXUSaQs9m/aUurTvJrX8vEPel/r6PWB5muBAx85OjZlECUzFLia4Ak9NJMFUAFv
UhtGTqXZaxk3bL+58EA5Ik6yjQjll8BUYQMLSw4tPtvRVDvS5pdnCxUa6phw9aN0MeBkuU8FC0kZ
gkuzCNCbEaOtOSkPxPoHYtcj/fHXJ+uV0PTwSLDd5qX5pB2aT1IVBx7dJRGGMtNMvUjObcM6g4Un
2fFFh7Wt27/yk0RXxHiHmzVNXLjrJqBYmnkwPUH8T2XbEPK6oFC1QCaNxV4yyhw5NzPylHDmca//
s+zdMez+bx9lGt2Sa5t0MpXkFNWUL3dBnSGG35GojbG6edHaBETtNa/aus+ETA5xFoC8ngFqkRku
c4huQyV9k+3Sf7bOhkYoFpEZRkgu2o9d9kSkZ/HczwFq8HvnWep3lCbrtZBJ0UtKXPT9ngPrRKeI
VMi3H/mffe8J38SrqMyA6dp6zXdUKMQ0nGs77E5xYZp8x7Ud8v537trxtK+y+TeOVCgn3E0LDhKN
Wl0F61Gn31ni2Qc7l+Tk9VlBnADXQzZ5/MmR/8zzIPW55UZpzDMZuEiHkoCMFtTDvgMkqMscJs6a
97HoT6TkIZX9EB+4eMVSpqa5dstUt9sDREgeK35iWbOsjrz2HxVzgaklaHxJeusci5TrxjecYOt8
AZmsRYKqLyKJ9APJScUod2I91d2oLf4fr7L2SsuuX94LnNgUbXcHrpEA+aQb7IlQVOXhclaQ7gtM
RRhpBG/Yez47usJS/c3DwGW/+0au9jLyB9q6mZ1KmOFAWYRWgkR0WUMv1FHz7KVIiUqdBNEmQdf8
4NzL0iL1JPLpsXo1gD4fzP5pxGUxPUcLT3gTdZHRRNNqPul44qa/4MA+CytXifqrGaxn0ROj5Y3C
DG8RbfZzlAFoZtebePvSEmZIU6+yWM1tGEnX7uc+vzypUnkZ2vWtH2KftWcQKaJU1XNFtyjBzG2v
aZ2pVL2Q6U10wRsYwqLQQU6+LeboEtDAo68YF6sxXTo086d7SsgDx3IQeTIrvGzOtBEfi2U4vi1b
NVJEqp4+O2deEdpsjpZG1lVNoLx0C+ipB+3w9JlS1CG8XDmwdBvLQXm+Dx/aDFaZNIEMwujcicDR
ZiXoV+/bBA0Ls0lHQ8ADXRuFDrVJGmBEPHqPQVgGNSPVK06LInG1D518dGEJG+JSilqczvIK1fIz
ebo2P0MKe32uWOWzvU9Krdi4ppkrewzrrCSaDn5CWvhDy3opQT1610P9IvHO0544YJr7l05FyNtG
ThtczlVpaaPGIeo+H6YFR+PnOHR9UikXOsscFr7o30cy5y3N2C9VAQXaWENCXol/YwDLRRTxeZdb
Zk8CS8LiIDAEWFpiq3tj4WpJcEvmGlfWY5HnchyD9bRedJjQwF2BdwRA3khTD+ddoYRZYzA9ZJbk
2tXHu0k/2XW4MiioWPBB/VOjrLOKIRuhaUEl9bZ8l+BkTyrs5qyS7p7KuWnulNxAYnkIuziDPjqZ
TWeD+bVdb2JBZ9jFTw80eLNjTNwicBcvXt9t1SPZPY+8xoQcUifFkHpvrfM+aBLttObGG4y/W+/b
2OEG1q1u5FEWgdQMYgzxcMFZJvYpCG5uMgYdlKZcrLArRZftGqIT+S9XNBAFBb5V4GBpl+BiQWG5
C5B1q0mehwNgVkQIhsl04Ram5itCU94Gl6vhkFYkYW+giRtZr3Bg4nAJhshTR02NOMzdwSD6cy9y
FU/LhUFP6ewB6mo83QhqF483fPwkxVNx/oF3nQEteilWtL74uLKxLv0L9evQoTkLNAOx7pKNG1A2
EruBU0oEaHL4SYRxiizS4p6lqTW+uj03cm/lEYeQKxKEbOfAeLJjDGKhwDtSAKxLAOh4HNcg6c4O
9YRIXRwmeCK07xqz891CWAdpPNZ5+4k5Ddcd0VFU8YY6D4x5URwEJaevfdlTuWMJM2X1YBj+q1KQ
T4WvHN4+13J5KgvmXI9BZoufLkSf/GPjyOFDO/6CZ8iymdUfRc90TCLxpKznPind/4MuBb+UUmyJ
yfDu7YVKwK4Vgd3FIeK7ZD2nqmw0f2VagWfD37MREc8cdX8313xdC/TzK9FJLVHfbtLENQekR2r1
zJKWZA8Q8o7EbgUQDNzE59cnalaEa7GfFNGSSsuK4pJnDh7+emHKZMuxHb4j/x3KbjC2DsqtP1em
quuV8Dastb42k71dKK8KP+6Hnbddf84GtKhhSFCgc4B2++2LZglJidvnNJu9xArP4lbMElt/vwri
hcyxgEGwn6qqNVkys5XiwJjFhRBTtEFERZN7HOrYxSZ9y9IxXMPOJaoG94kBeaB39YyrpvKU3nSM
Kd2OE+gue9G7SXD+wtNe3uvUVvz90HTd5HEbwk0Pcc7p8xsFpfJM9EZxIwKkmP6lw/CjUL+qhK47
XFxuc3Nj9Eg3DA7kmtQ8cMH50bKlPOdCWfUeJpV9kxrsXbygYEt4AEgVO6fIdMw5dENKUjEdQPBz
oaVMs/n4/6onOFiiteXfsrB8yxSFhzaQdWJSUolmkoilaZhuL+KLDl9WhNilGNEGGVSHbQM3cJaL
WzmvH+RW8kC8TCBSbIGwrFL7Qi2iSGvWb2aCnxj6hnmecTKGmxgVhtdv93M3jMekl+DE6ZVccO3K
kqEWaCvzlnseNig/NSKkWxjh6Ggr96TCk1H/5NB6iW57w1kL+HGp2v8492hvKWHp9njHGdSJ1OUI
G9t8OSnGEksSzQYqz9vjWQv77bhAwLQfILPnHL+UkyP8lnMvP6QTdIKboBm8DSA8JLXaIIQCUyrx
aAalHei9lVhwHPUAgG21Sa/45nePUQsBhVGEwfesSpcLIu3hi0nAkfmJVdr25qcZCJoNk9n55sNY
shhBls6zQ++ZUSA+KdjnQG57YY3aqMOlr0GQnLZnGObW371zJ23Dv2tnmm1XAOP4eI334HCKHnwb
Ss4BQVOZadsQbmj0B0d0f7oHBhDgydFpWmlcytulR7IrABX942WjfaB5PHX6ND+s8aRDEY5Me7A5
kTAprwHK2KwkK4QBwpyHClHOhGTAa+90jFu2M4fgAs5OLyb7Ska3vu1pUhCEIn3i2H8Db34K1plU
+KERlFFNA8MjaGv6pmeqIorydhFd7dGvxdEc6E7wvrZlLis9tCKKrKx8xintOrGCDNRU5fmBi04p
Z9rQ56Uf7pmtqsJbjWWVVD0p9SVRf1bdAp3Zqmyk+Pvq23lGZ24TVqMIWKLpL6b7E5Yt8FFQftgm
/ds4AU4fshdPlRtKiNEWWKJ2fat2kexl6YfnKP+cVEh/CfzpOjxBctlsZOC/flD44C6AIkGkHRw7
wC2c5MenuAKxEGCbZwZKUm84UZbInG5r6IkZLsELFkit9Z/PjETBjCnm/7gnHKKAow3fm2BX0YGE
3c+ZKT9GDLSJrX9CD8q5RaM/j/H0wRLvMM9vv554f3b3SLhVvzUB+YMg7FiQ/aaA5HDWc6vq5ecN
O9GNlRNmeTatZtzU6B+1czD82S8U5ejwBvbUxIRxj7cbSiUVZjexA+X/at0UN+3N+9+vUc4h2XpN
uXZkcjUfbuAx6PMCohzUyQgmVqbjSO/xNzepvez19UyB6rgDlX/xvw6C2mhzThmhuZygE3rW6tO8
YLxER9QiRAuDR9/T7uoZ2h6VAT5nK0sUTz+9gbEdQbTN6YiY3bODYGrYh6rn6svd0C5k24dDRCId
uDtan2779p97NOrk8v99GqAeDaCKDu47zC+NikvsqZVxeIaV7I3+JDNp1ENRfyV5kromJykNBblq
r23w46VeTA7fEnADINYmY/RVlkVWy9JT0OajDPnMht+3M+HMGirdZCnVAOuKRahM0okYKrTZyf0/
wPULVjQme6fhLknnxPS3yH7AfKVDRqzuMdrEqobpJPRSpEZkYc81zP+QAWvXDwCArKVp5ogl6k5o
AHiGSP1+8BXK1Kg3KcxK3x77XucYTcBWc9izyf3YciwUEgbzPy5hoy9DEo0i7MWgSrsJUIPxKUu7
0TrNTMNd+7w1jrrJE0NAwy66N0W7VhcuPRnqChZ4YiYpy03351/kCa8t6AHI2xsXUgI9M28uml1F
6OBm9Tv5ap1jSQiVaM3tzCW4LdzdoaYbAeRCwQvJm2zDGcDLt0EVqWje1BcvJA46BWxlodd0g2qj
Gb6byOyujTgxZofcJ8DFQiCeppdvKFctgE4WTtJl12SsXsCbI2wH5EGBoPK5QAgQwUL+0NvwOg0F
VeBqxm7smOtE/9S6zfsvJI+D4HKbvueoikj44HtgSI8YvzmUk8bhLfjEvD12mX13vKYLBdjgdECc
O97r9EGXMbD8m36s3K++MnbYgHrOfuo13rOn+Zt15XSUtQwitzrg5TPTRmpCS585W9EHHfWabgoP
V85AOBe5ZKhYsk9BBvbCqiXnKhQDj91XuoWWVcVRB9kiyYqf4feT6TkHSyC8U9ZYkI88YvkE4tEM
FwKujAs7TFb1n0JmSJf1mS5zFFv/Ppv1jCserdwMW+ALlx7YKpbkUraHtswk1JktCg8GZHrFFnEE
NaWbxl0i/hIA87SmAsteosQHxpJkGliXaUCejD9Wjt86aABsoRlIbYo7Hw2+OOVdpvA7J8eWInt1
O6uTuC7tDAsLT9guFEyos3H7343rvfeh9CBFhi//XYKnwrZ9+uRM4Z1rqcPTyNM1Tehnh8fpkckj
AczNQvqsatFs5CXbwpvAemOsn3BUwAAMBJMev7XTOsUnCZgR/MPYmjb3K2lDg3Y7WpBkyqz6E4iS
OjT4ErOSwc9VRtPuJAAvRiWwYYH6cHm9IQgctH3YrDP/E3Llk5e6rlKkDtYjmxZPKHBW9pCKVYTM
L2jzBX3nqqqfNyg+cDQaDhZ/tmEM8hujn+05mntcscTagVC4+FGh6/wvpZw7F16mMrXUbOksxekq
4sQvSnrq7uKGEx/NWAXjGImktuiZdRLBYix+E6WskApZDVWl7KsDUeg8aWLKobrEgNMG5aOobUXt
n9ouIuk/cHcnJKiCfaXZxJWMCKNnhjzzEMs9BKVl/9rtFhZKXmu2JvRGMKxPGekSzeCLreUM1t8w
s+CWMfuwjdNQGqN573OSuJDznWWXpxANYJEKBhE3pWIIRloFoGVRnAwQ+TT/XYAZRiZIYYEpHZrX
Y4pyCM38rcNnClUJx+V5xnRhPPcmH040KVBKhl3YlxraFIuNgFUGRnL7Ydp3jCzkNqRGZ1jsojM7
u1G2ZV295ozQvnJh23gb4+Xn8gmAoJCYixMTv5IOgXJAwuTbewxifqX4FK+qovOhJY57wdtSIoWH
j0fiOh1/6MzDr3pYoM1krYnW7QhjDIvwI2LlopGcxDYoGr9GPqc+g5e7Z1KFzvzJOkqREj38SGwp
/3fF/qP+GVrwGaI7bsR4UqzwS5hpydze9VuLn15pfPlc+IAnyvuXxuXlbHN5Cy/SbNTGWpVyiqUl
sSoK60SyibhR8uwrpxgEUg+QKZNs/3dQ97SDHCF/T0HnShTbdnUNImtGfwSq9Ezblp8qNJJmeV5m
B4JTlwd1J69nnhFWMNZms+wafX6LsUuv867uo2r4PAIeQIUjqmREYaBCpuLNiBunGJrzVfr67UUa
vB2ZlOq5Q0ZpJpaTuweLmRSO1a7okq+1X/kbxKEEqzKQ2f3zYZxWtMehXuMvijU8QKOSshQBJTfQ
aDYDN+cZLqyAvqc9YUpOu821Pv0aYnAp07b8sdyCcJu4hRUcdZDWfr6bQ2v2YiVKv+/LIAVfC3xG
4v4Y4OU3aiS0SkRBaM67oHvSZyJB+Eb0ysp2OpZF9+Ee6PbnE4aPMLPXlb8bvkItBEH0Wbhfm0rz
tFuAYlnY+Pgzlxg+ls2FJ4UbM1dvdwF1J7nVPrsraiz+5R0AlPNdCS935JgMrdb93RiCWWXr6FVg
8Te8PDDa13GuEH0RZtU+0gKuFg0FDLoyAtTpV37Ph1cPbHSJKd333FOzp534NO8plq6vhPcnLNds
OHHUFTvHV9FeNkSmwzAVFqBO97PdB01asZgYsXF8XMZ9L35fSykB+luRYB6dNjC2gH5LLi6nFtXT
ztjMsO35e6ZcfPBDbxrNavodZF9HIixeqkGyPnbZ63/d2cyxVQdLKleDVhvdlv94lB1ad0Gfp4pB
Vpl77jF2KCoersUa3i7iFtqPwD87otjko3iYqFg+x43CLfpQwvNDWpjhh01bLPkLZ78MOFZv+8FX
OLBAMrzoBEFX80z9PsYvtXL34mTUvthAmLn9i60uGhG7t54yy9D7GTIdwTYHyJPkcYDiEPskPz2L
LCuVqnaM3m9OtiWCXJ3lv3kt45h1x1eY3E3wllEbbUVWsnF2RZMFGHvHnz3q/CAqaWZ4ip6oEvSH
x1KRgazNKiUiHpLXQ1PzQv1Bsji+OzNsSaJLbQLSdKF6m60UTyJF3hfGmfE/joKzr1iLD+LMw4hB
zAP607NKsXZv6grPNE7BoUHJtJ7bMQip8T0QBwIFVVZRVup8ZCCRbuukqfYaS/W9rACYXsa1pvzw
cmQeDdI5+Rf4M7mMB7FVEyLlK93GpddS+I1FndwjlfZcq00NehtccPD83RKBVhmj/PqYXpQrmZ3c
ndqLck4k0/oep/jrBqTDUI047Lfgb4nkoZJQJWdYo5eam92ejM4K9Muig8TErPX+URe0yRwuQs5r
Olxvr/di1VxzauQbaqa2SKjn90ssEgWv5V7ChdJv/rdKIkqcv42Bk1X0/8Y1wNxOAsY6GbO/kVDk
bVrVE5wvjhfKLJ8P+Z23KdXuruvgq9rVBfIzI+CEn38Mgja8G/aTkC+8w5nffa9FFARlOa6rYyC9
yGcWpcSMlbG9lW/n+VPW1qJ9vNAYSNZKWQDvdGZExQ/JffatY282BuqxInV+In3Ulyj2Cqnkx+lo
a+6q009Ea1Qie4R1VbaYffjqsCOegTzDFJKfsRQ/7nH1aGwxME7VqAke5K6WHBD2CkRwURCNXqsB
dvridJpov5DC6UvSTMm1amrDW+vIROdZlIQivqUDJaQ95fFpbK2wSWQZwgy86z8eJPhUgU9OseTW
BTQd3u6CbSalWlX8J7+++QbBYfHgK2RGqE7yT14MeSEBpAHk0536011L6oItRzfH4kxBO8sdyNcx
tmxK7rKATCwyimQ3ZUer5vzoX5G4LmkLOA5/T9eankB5aK4zIpjsPniapAs+LWqoqeq0prxk+/No
uF0huXYxD8KWaI7QdlqzxR4Obno4bEsYn9FZvPvu5fZMv9JirPG8wt3FQJgY08o+XOL4ZtrAuzSV
5q56MyzKqcaCzkGVilcBcPYpdXWX76IbTsDzSXXleAI1KRXru/7Q4E3U/9zRnhw9yiuxSuyBo7D7
dgXQ10RIxRovbax88QYGqYtf48E8bIKyakwdIP4SLxLmlR/dXuyWNrHOHqz3Fq1hzb/jvhW3X7GM
tENGAPtW4qxQ1rJUYh3YMn2ZBNOg1t5KTH/poASg8w7RRQTitEVceB8yEyLbkzZhbHZHHy4ydcAK
XhN03flpIJi0OAtB8qGuwE9LDNjrt+Hkaag8Nc83FPDXVIy74mkiBvoYZ5opv5jb6LhCneOWaEwI
BeqQDNv3uJLKWB0wSnNra2Iu8fC7UiVzUon5rZhl7dYMEYxxJzw5+XI48/X3QiAA7RO1ACoRoBzy
URpADpgG/aXt04RO//m3nK5i1uRriwhpmPdirJ+wkwMN+6SOynwu1rl1uKJeUm0Hqw8VJ2bhNUlT
8mgmThbVAYo2OS6UkYWF5up3HpDD+BYz7CGXvFD+TRqZ8A3Q9j76uLHodcvVdqoPyORq+fBhO+t4
CGUbWbwfPGWJeWwB5QceWaNrjGhipKIYndDMn3ZyQPQRP5rbStAHGfH+9kAfeWnZ1C60jJv4i5Jy
LUgtf2pIwBk56UmVjlhU0xHtekCCKf58pKMsRYriuYKEt9d/OJ+PexzFZXlm1etNmlmxSeRg+JEH
zr689Ykf8j6nSXG457hi7C2y4xQUZxfwLwxYCSu4OUN6E0Lyo6etWsJpvUeC4r4kw7i5P8aedt6+
KLc0kjQubU6bticZj/v4eteVDPFr1gwxl0YW29MDWtT9KGg1v+4Dzue+wEKFb8Dr99uPsSkYS7d5
sbwf0SkK+v3FUOqjgKGLqXOXc0zavpo9AH/Lvx8Y7redHkyC3IsrtHUg6NU+eBEnaIDx31/EqfdT
jhrtMWj85HAVmVEsATDt9hau6uIbOQWEX9CL6R2IzJRaMvBa3H1FNIcdYuEAZE65RN2uL7LXLOga
qzSgxhKVYG6t3yluTCqS4DqoYjFTL9B/Cf+2xAjPqEYYZ7p+lw3Dvk5uvvWoPDjfO1A3LsKq5NE0
DY7MmCE3Qo4vrNGrzx0yOZAT92JmmYrfPaav71LX1jcLNb6ux9LyNGzQCPNyFIgo0MzhV00/LRUE
2FFxo1r2axdBI4zWXu2k6gp4VxWBH630C81fwDs+Tas7nfEODxMakkQktjhBtGSZ4TAolCOqKFSm
2wFm6cxphV9iYTPYb46Hn2VpSYsGi6qRGwxM5+Cg20kFyprUpoMvKEVddWHpxESCEGsGXeqKlD3r
Nt/g7H7ofCzvIcaBMR0Z2X5eooofuJgtzF1dYjYDo72cyxisVQ/8OxP6lZJvrgFWrcoYCKCUOFK9
OJMKLm0WbBWrwzvuPwd33dSod9rEj9CBJU5gwCOp7acGLnhKKzF6EoL/Z8doZwhI0z8cG+JiwkyG
ygdfITGEYOPm+ZZe6xZHnFqYKZH9d75bidH6UE9WWbTHWOIipgRfKuX0eB+sP4Ciee6eHx3k6kmX
84HJjREVM/rye6v8Luh70XvZ6AWUaga0I6dsK++tIwoxQ24RQGpGqPyXe8RKJaKHZ3pqQ/ywhjrS
u/KCOCb6uX14XGocORWIXFnjIH5rANwsWRJF1KfbG/lEVGPbwPnUBh/2OBRaKCePTlxHj1UzGQvW
I+ROvj/vLRX7ss0TIpvsTA/xT+VCZObgJLpbPTHNOd+NoyPkkIXMDW1BZAXAmtj8A4Qitfd8JRVQ
EAnz5HXRJNFzwBVTSGymZLkcpgf46xe3J7imqC8olO7Z0P6Eu3GQ+xyEa760EYYLAfZNbpIES+eB
R5w3aY4HkghXTycFaoPiLMAp9iBxgk+4pEEBRY1JQFLrBrdDKBArGe9EjaUAYnwQyd6FVZK74X3o
xiZW0RegScbpANwcBmTwRYarD63fbJrcy+SNyrI3KegAMWYvWznhIgatR+DjLNyo9mKEHgmqgLqN
87ybUGGya1BkZfNeHBSy9fULPlxgXk323VgyD2n7i1KL63wz0qnU+UjIpk7Y6K+VLNJaZsBiXz3J
sNJy2XJrcqRsI6hN01hqmMc0m+XVJ4+favNAwXz8R4z/kHXxf+saaXYaSVBq9q6nz5Ouu6tsJxiI
5bA9syHUlDQyjEeP7oRoJLVjepjToHx89PHg/OGss58eOKWQCJ+BtaSREPU96vWcn0ZPpvT/uXyE
muekIoaT1SxZSe5wvZwpH0QyPNQ+bk0MpUU4E4xSxBr2ZMl8ZtTFT8eZZEdrAImfoFiPNwYZ7Wwy
2ZpOQUmH0GvWH3HfnICafSre0r6jlYc7XPXLjQck4Y9BHKGbQkwcwQW1QmMb4sVmLwZouhVdHLel
tJMKpx6Anr0BKbg/+OajZRXKl+tW8xxerUJNpozUTG2wlenESc/vgaRUS0P1mKEDbM87qmiPZH5B
1ptuPmXry81osXOYptA2NqGuMluz2PS+0IozvnoNAlKu41qLoPAilfiEF/qwLPxPKe09kPspFrdG
68Y8gEdNR1BxCWGEi0hz7x22rUmDndOjhVqTfoAI7PasTqs9k7XErfMGE3Cctp2qm3etMTCLSNOO
XKAHuf0QKqndUsAffXTk+F38scYpasDD+hJ1JuFZuBJzMAzkzWzsNH6hyrb9KEGQKmvvlv/zz79R
mdEggJtRbOfvk7FlXuY1JuwTaWJhcY0NILD2iKbiX/vW1gIej/0ISexWsslgdeFBTAT6tfuCUx2O
PnvAHj6skrtpTwuvLSkFTknXxlBU9V9PVZk34a9TH14gDg7F2dcpRZX98YAl5+DJmAlDc8p+1Ig6
ZFEhNam+UU+d9v+VXK5TqCIMzextl/HOd8Qe0mCCAT/+chjgl87pWQiPlEDVVhMlWURdgXADj/vB
QQoyMg0w3+fW59jilxWG8jpVZOBgVanM1aZ1gQUN7xUXMJRfLtV832AmymYrDWQuYqrhaKxePBl0
3U7pbhVce6jkgLgNM+D6aonDkDs+EfTMpqW/JBt9ZB1ZeFyP0msE1KmdSbdl4YB3oMwiyK2o7WjV
pZaM4YrP18vhkzZSpb+olv2n/N8i4erOXn/qB1svzJBbiLM55FxHesLSKsh0P1XrgBUwOWcdOJhy
S2ZZeReQCeJtHVCe/PGpVi2QTR4XhLxVzmPicTUVdehuuhZe7xP69Tq7+59YMcUnOL+pKTXwGk0q
pTp5oZibXrVA4rRI1EnT81L3VBR8Gn1k59tIpU3uARoSb8ylIFhBvPMZiedRGdqtrkC6qIlah62i
Dai3WbzJ3ZQAvqFIkd1DxFT0b3JtEKSjKjAuj8FXBP6LJznWQzRH7md3z5btnn4da0yGweLX1QdX
iB9oNPskOBLDQhh+MuT4VMnjh3G3/SegiN7MSL5pM2ZFW9jYPGLZ+hs52otre4lC9Ad3TxNeNpJZ
zMNaOwD+9McWg+ARL/L0EIXQeMPmj56h+ISHwlHwRWO8UWymdZTO5an+IZxnm1dK2gbdVsN2F17I
rx9OdStq2+sl28xKmuxY4dAl3sLQ7oNAbyEiZ3N/20oSLpNzDbkma1po/Hf4GT3e996gtn7I60Im
WJ4Kt71iMavKKWjiv+D7KShG7wNNTxqwn9j4sreYFjvmHlfMci5ceyBCxI7QGXK7pLF5+359Fri5
gGTwCXkugZYdFMa5OUQ9ilPFA1BV5eGEn2s75/8gFCfDnuznlJi1H8H2wdYlgiUU2g1Mtx39U6je
3062f1BXb6QRpZJiPuk42b97nzzYFfis1o35avwsk0NT907Hh9SW9nBG8nonBZsJA1jEUYUEdRsF
XDrLFfscRxoZD3OPD0aDGM39EO2vuOH7U2A1q/Ug+gaiJkMJGMUZb0kbKzaTuJY6K6AeZNTi7WaI
5MdFyvJ08JBG8JGJBbNU3xkz1DwYmAUIDCyE1o4yM+ex0B+2Hcmw5jA7XAhj/KgUkXc90Jmr2W68
zM3wx9BxwrL/Mi7XARL0ehETGq/QZC0CWl7FRF6N4IyzXG4bPBkL5eM9KeTzDFP/MY3As9aZxsrr
Z44VJ3cIJeBmra6Kco2hjbtaWp+qU7KXPpzYN4Aba4FQsxQwclrkrsbV+MTmN9QoLrZwIEyQCQzz
l8msXApXSL0N7GaZ+9I/i0T/bGeoVUOZGyfwZTZTItMXv+DEoiMEIaoyCHFLBpuRcQjZ77dA/BWE
v5+jU/QnyjJRQGTxeo5LvMcTXdrsN5Gom2SnlT1oTeMslA1nXFmXnlwXgvI4pjkH9mPXOK/FpLNo
Q1fmA1ZBJ6drg3BeDZ+btfcpAmNGy8xzhBlRqZS+xiz4FkWtXKMm8+B4rP8HbNkozNDywke6xgjA
n1Fn2VUa6I24HNMeHxUfNvpVhTqHgcKTwXXOnf0uhOk8z05JVrOcwB8BMrrXM9RPXVpth1y5ZvvN
u5bCYSJIgQmttX/RGE1Kzq/jGA42Sg1dEkWecmyj6jiIAVVPA3sFUP/i59BEmYFBvLxlgDg4GXSw
r6deORMA4zlFkGccQE6Tg3Xpv/mylBmfYS+y1YZgRLa1NDHtMcf9oaI8zccTJDpoWPKBYlWNZVLm
0XwwCXz3dV9vLRafw39jv6hicbx7xB99SEeGNegcwwZxhhfFu6R/Rmf7wkIu0V4/ug4Ce8pVkw0O
gdFPlzLq39pL5xa3AcPXaklKXXAMFgltpIewXtTtZzmdlvlsJ5Z7YvSYxo/qLwNncOXYWcLQgBwQ
qAbIb5aiFM/PvS0FR8UMS21bdnAzaWiA4MXKfnSbKcALNW7voM8VudP0Vc4nyftQqkW+BFjLkvHi
KJnBnrcDjlZBAm2ke/ITYbeN2kgXw+K2E83Gr/90roY6eONTVjejV+IaU5h9r0OsivHa5m9mgwCa
vUBEo8WE8b26yB0irSVVlu268FqGF5NGb6zs8ltrnK6HQKb+PUBa2DXCglDiV58AzSA1qufG3sUz
bfQPS4L/C1QWYgJ8ELvlxCPMW+H3+zD224ioCoD8KIHwjBXbu6h9CZeS1j3B63BJSZre9/3PCLYa
/AYmhB294Ss3TKSKv7kIFlEm6JMUqoKyD65Snd++X4PRdkr0X6dPiGE8sXrz4Sn61+WNEzgNCbkf
9/HzLrSSgeEl7GFXRlc6plAqgqsKs+fdY7/sPgPkWV3boKrgndpwJlydD8mNUH3J1V/Ds1mvVn4H
+5aFSeqMM2p8mgPO2p8MxBQJCPsz/tZOgPl+JFE1YyP/xn4wRsTchmj5HML2lLCvUzPt6/4nanne
musQA3+YWEhYd7A4mjknmiy5Aj3iba1dyndlDjuJldjxytLu5P8LJZTfsz0BGUERtbwLz/d2Ijuk
Ibo4A92ZGpCOLgh443AO3QrbQIDupnO8OkdayXKqretTOtoma0znkfTyCQ1ZlxwohWcWP8CB63F+
a18ZCFLEXB5e3Sj8JOIpNi1VzpDnmKA6NYUBura4mMCcsqnipxY41P4AF7wUriKTQRRVxLEHW4x0
mdlrOVbXpU55erC+5QZ0MEE1sbkdxgI0R5GXag2pIOzWi0K8WnRG60kqc70EXA2KjeXgdOfCdp7V
yXbYhAmRWrLxdH4FvUx3tmx/InAmznlys6gRHMVLyg9weTvYbwCjM6NPgRfPMHDztf8U8L1rtNsq
g5iaLdce4ky/mUgGZqMB8RmC/l/+44B22HvDdh5Re4nOb2klviGHpEfLOrNsD2ZTaxNOQYOFmJJ/
lCeXhJFStZ/kGyq19L7sLfVn3lmwFHsy0Fap8bvyuKbb4hXpAc5XQ91BQbvDTyqUEuRqQwoF6FtJ
XHSJZdLNStF1CJxrH8iGU76amtDPBaruZ/6O0CNIVEvWzSmiHR7b534IWQKQEob7fho15y3RZo8K
F625thZd3jf/RrHnr87U9ANn/+wFXHY4ee5LB/eKxZ8sCWRpPnugRjGEt1nIv++D4RbsgPAMO8Mm
ZkzIy6oaJfRkQWg8/IJQAC0RtlPlhMHE3MvlgWWqbtPDIQcg7ApTYd0YUaqw0gNC5/Dhfz5NaQ/0
/AlB0DX3s9rumNVL0nSyZGLn9Xud1h8ZD9KlEw32Bc72Vq8303Y323Y7X5GDD/0S/6qAuWYkRdov
1V6/9DvTEANtet/nOJCX5xEgjhth1+oc/fNN8dkIC2GNpqrZQLn7Jh6vYCPQLbFUrYtqG1Tsr1Y1
7UHpbP3ox9Y+oRD/uiSOHT7l+uvV/FhS8f6UK/v0hoFXXKocvxj9vVeGry6N8mOsvS/8vavac7zT
tJK+EGqncvx0KUIooy4GnBm1x5J74oW5vD5mZbIYK3DXIBK/LIhWn4niMN9jFkH2YopZ1yLl/PN/
NWiaJDSHaafyQJN8rjzrQAUXUZ15uNbxR5MgplFL5md5OBdjJ5horan0gQhy7PHW3ULSPf7NPlVk
fNSnB/fj/7poG7wdGD6Zj7f/72fCUXA1hjNxGi5mA3k92FRhRfUp0QsUDRSaUgy/s++hK5MdwHw8
vCoOZURnQcClFG1vmHOQBOIaWgyYFEIDiKzEsKNa/x+4B71114WUDDbOzsqrASOhiFBzPOciQda0
aYSbb7xM3AUm7k8KuZ+Io9bYyN+vVfIIt652ioMclQjkZ3GXwVGRTud7I7piFD8qhMMlX0W/7zNn
iT43SDTM6oECbC3wQcBUCXEj4SdAlI+0XLGH3NhPn6vxOPxJFBrWYK/90dpsVtW4xqFtID+C97/z
E1r36kb4DFCKIWk+sH7BiIyCMHay7PDMPoitM3po0PofZLnjJ8f2/6kW8Z6tIT+RXMBZBv7cqHXa
41N99hCwLFlUK9KTw02mSZtj64Oq4+zUqIZ+wqV/UOvBV2qQ8j+CgVCjM53n2Th7CADTrYtvpvdg
0ebTIMFBRD3l7+I0Wk6hhxoZ5evLVplUR4mjmkIbe74M9v7pDxA0LMx39xHpZNc5O6qtwhhaQK7M
MeyjCgAFIs7+qombd99DUAc3funNt+AE/qUv/vzdCnrXnxizBk8tA3M0uimqBoQGbSZMs/vODbLq
gkvXOaUy+D5tT1tiCHRMSdjjG99lUMQBkxT+WhJvOyajxap3+96Wi7YKDfAx05/AaisJTknv33eL
fip+05AS0Bd7oU2q8CUUt0sufBkV5LXeYl7PKMgBtON3+2gVh02aG0v8PywVROyJ+S9wrSDVnDxn
nIkL5iX2CWSkFs6jkwrGk20P/1pGhiTIr3DGG6Hp8m5W0aZ/PQQfl5oL1lrEOptNyj+X28yGmxHF
y+1jXqRmdbJQN2QeXDocZuBwn4FT7tXrEGhjXA+DsMkltiWxB9CVE/kg+qnMQgX5cAuM/PXoxKr+
2u/TMtEjWr2qifOVsCy6t2HJgYks5/TGONFs//pLMXsIE8gO0ISFkbbkqzc8L9rGIisKcPaPQEU/
o87drCXCJ/TFVPPyyxONrWqes2cP3CTHlxTy6vV/NgotkpLeFgrZHze4lkoO9uhuXhJWvzuqedWL
57klww8dWkduye8gzDoHpM4A+I7Jzv8dlO7NyvR2iwNHN6wK4LcGSW0rCi8L81p88dApNZlYZvAO
V4g49cUt/Vc7sgAWp/4J9HoXmIuafhAbeu6hstPNeNRRow88//rrWnC1VYcPIKunszBQj4WDWSfu
PiBEpvhos+bFKcwUvrr7OPfk+0qat5jpP/Ef1ZvwVonhXzbAwWjg6+ryUJ6a+kpbJvH10gFdejt1
P7q1X92w+sSFPvpVQoSz42UrtXn4/ldwvMRHRg114WfmjkA4W9ITndr2EUI4WpZ0QflS+0f1e+OF
N+/dTirfGTu0g8U88IE/lunAFujeVXCmcezisihPC0ZfGQ2voPgASHIn34UOD76YyOW/uieV/rRs
w0NUc8zpHgDUINfzUOrw9hjT0QBvZnMUFR8iGQj3NMbLNPz6J6wsBWAP/b3LBj1LqI8U1TbHCPIs
ypp/L7f1tMZl4WKAf6Lr/NtBf2mmY1/WOiVJjlPUXmBG0WWoCJRhhMJbtb1vV6AffBLbdlZ06eLh
jBA/3MH2UwJKXqnGJFZqa2CFSVet1j585W+bpZHCxW/GtwTGdz10aYX2gRZP5yhApZAhHAEeu7Rd
QLXsUsz5VBfISMi98nmM3sfoFderMKg186PR9RGwKqy0d1oxcJK+zDeJPsx70zvjuIjttXooxIoM
Ttf+3lnup/cmk1RpG0/x3RLaC3keNBuoQ5MaeiRfJZEVyRmLWA0Vof8HWRfQ3/LfaCQygMf9x1hd
ml5JxD7szQ8F44jXn2Qf8efhXj0QeFPli6052xRwnSzX1IEFnJkh6DL5ETWL8Ay47Fkb1aUDelNf
yjqsOUxYAQg8aDNQqwrLQmmrkTCcholqSsBBL78oRXfds3HtqPPnVcEVReMCDyT959V3iK71w9qk
6fIzeDv8c/9/S84kpCdK9tv0aKGo4Wl/BXf8D7OSoe+sMzT7Ksg7QDzkg3snvPx4RoZymXSCXy3l
WtkmSCAUX8ZSfU+fwq1muizm7xU7vKO+PbGEbPknNLxFB+6CysTLneQWM4o82wJwQMiZqZgIzFlS
Kbb/aymACxCcnn1rRF7nz2V8eRQLlW+0dNDfvz94Lr5R7HDzI2IqCbFe77gqeeWMwrQIUWPyhGgq
FPa93lS+QQnLfjlH76soMdYmDsutXx2RBkddrifYBgZmaSoIXA/5//EjIYnK20KOfswdTylpM67O
TUKkoi/cNxyWS5TRzPA13SaZfgHwg6qDC4D0qqnmqpOc69qAcNl2ZlwZlL/NbR3humyAlkaIwkEI
z/Yw81IdrPR63lEdIlz99dUAMBhSaUZwME7nMBb5TKG39SJTiyZQV7VLVQ9I3NraU1PUr0GTJwpJ
NRv3hF5KoAvbEm7KWCEe1YZAx2WSMzkRVfWMp5nGkF7TZmevXMrs4xci3P0u++6CAR+UwmgrIBBd
7xql23S1oVYG+6nPe5fyjzvYGmB9iw02DReNoVMKRMVSXoKni8gDvx/Ze1SO3T5CZE46ZP1oHDtL
1JN0EvVpkCqgMfIPs0S2Olhif9hCpBeQaEMyIr6alxkC8hiWMOJMF/IA4Mit/vF1Yn76gq+WTO29
udKBlY8Olu966KobTcpqpjHOyM//nPwy/ZQcHhZ/yOEcjMQA4mF4qYkJ+9s1u0sUWU0zZ2ypFwNH
cLjsoKhwyW99WK5kIdGAZt9vfXUALgt+Q6bpbO8XkjL5zbcAw4HK0ZLQ3oM2rVQD5etOfpN1Z0gI
pLue44N8702KKxFMJSDQYj5Uonfw4/0Cs4loZNKbG+Lmg4ro3P2EwDYF9RreRKDboNQ1VYVxooyY
FHS/PQy/bH6QFvU3QbvyhghvuEWziPzu/MpLRjIPEmH3u0TbEOuMo2184oEco2qFs2Ea5NwB+ehq
OncIzNQAosPQ+txpXexOMNMpqKODUatxVwzqiwLDpd+fke7KdQOT4kl5tFrgUaDzG8tIFj+UZgwR
wykF3EB2de6tFBVm1Z9Z+Csf/13JLWK3vKFd9IGAHNJqlKdrOJ8PyVPfY5DmoJ2rdXrHsRl1zB9k
v485pnK21e+8tjmyi19U0lcC+cxdXMlKqLGkdbTOCFO5UwyFb/GykfzP73Wdh5kt9uM1ji+Jk2x2
he9lYOBtUoXbdHgnBF1jenR/ZzepAbl7j7BrxdXb02ZcHbwVaxldKz9OcAldMFFv5fQm+EfekENh
JtSk1T72Wb98uYzcI0Pkkzud8uN6VLGF3f+Oo3B6zkpSmPuOaU+uSUVLIJdeKUwnLmJU03Rfq3O+
MMthrhjc+Xy//bF7qJTFmfiPa3+Q7+Z5RQ9Dwy6BkbvRmY2q0hDZMlZ1sUTiB2bz6VKdSRmmpSww
haP4pyzY5+t8CSQj+CC22OX+1xkAzg/LbWgBP/VMKp8wSyHSaf8KOpvT1gjCHovANt4DiBEYsZSM
roY3C6+qnKaKgd/StRyIQdK1XUjraHuQL3vaWj9SCjI25BYJ/r3GAqcLFi9tJiqF4q5k/tm2P/Xi
KBG8Iosk9Q03zUlr2bBjgh9jXBF74kIr9iBqxa+8qL+we4LKN17wZAiYVJIXdjzMEDsaEScincVM
4bpIPLUcQUzl9nK+98KSmrbs0wdxVbaF5vnqVNEm8fL4KISJORUvnMIbEvwY7+Xm/yCXp56O63ca
aH/0JY/xuOwsxLietEHSfXvTFM/NcSqZPayrNHKvjO4wgYlJQK3qkkoHvSpwWng+ZL2dl9ASgVgf
yhzo5SgMpez9uAc8ONpzkmT8QwkLYRzuCvktC0zqbFSin2RY6YpsItMpdaBSiD0YzK0RgzokRw8U
P2WlfYSDkEvft5q1nJzA8xr6SMwGyR5WuzTQW/gEDX7+0MKm3Um20e8qEJFO+MzbrDzTwu/Y4Jcx
gvOxbxcy/E77g8F7s9eyD533FsO8MPioItLkHsYoXOjNkxq9MvIhP3ETJnzu8Ohrt0S0v6rwsbFj
lSAE3yPxufOSsmQD8t0l6qRw5XPqSa72rrXZ2oC6xSzgAHAhdkQkvQDGprvuvfJkw1e6vy8UlN/f
n3RpGISxoQU0qH+TxNxg/jsEUjNT9ePMOn7KDuK38z73YsiptN5NGAMn1dspJPmsBud6eYV98OSS
h6ydxEfv3xrgkEkOJwaZ4id0nPkrI2u/BFKLkSXCLM8bxnfHcZyaL4jx8YYvoOpRY2/4+0b5oFmN
QNhaegyAbsxTS0oeu6BgA4axWEIovibFZKPlqCvrmsJKUTENPrgIs8/Jlnekfn+d/bnQmbIbvAeA
qTVXPDVz/c6Kijz4GYkFnlD/7T/bGlXnaJi68m2Sa9OzVmMAm3ikCw34zLVWNlxzpdteWcuAun/q
QZ3g2ryj8n9MyRicjL4on6qTbipCARscEIp6YTN7gU7wJBkAEg5NkEjFk09hBNKXPX1nli6+ppui
/v8wEx7pYwzWqYSxt18fsq25pF1Dq10IJZn/Qp3rnxOSeJ/WFWtYg0dtbV5SOCXOVbGwFR5oxYhH
WFtVujyz2bfDjLEvrBF4bfv4IaNJhK2MzbaNLpx1pj6CbzHQG/OXnA2GeTbI8SjdpISfMDkXPCfk
3em2kWnkMUB5zhfDKpLzN87wkFsNds0Hh9O2gvE8Pa0F87on+xJ8BWZ3N4QygxVWztWPcIqxG5D9
NviGZO1f3VQi+TgovLwNFGnx33KzKNvr/hn1TA/Gw3DBUvmpU7FMKhTORjl0wscyrNDwzhIpgRSz
6TnpeBupZ3Jtdl1fBQrb9OauGw8typsilkGMJAt1PYiUt3/SKK5SH580NpciXeTYILuioqMh07Kl
sUKpyMYnU/n+w/fBqW4O3lqo8dAq4DYDMhb1DihOBPcEUIgpq7hcFpYlp/DgdZFjX3qe56hqFjQr
+UCuLaQCYi5ZzHVrNIVTU9gf5rEv0ukwhre+VPuNW0STSimQlIgvxklyBR2i6upAcGOGUw+c5nIr
kLDkWfjKO6D2tIUX8zpHLsW/HAvd27F4uh3LZZLZTVgBvc3Wv22tQCxWceAdtiGw9ntwmpMQLV8m
xS1gFTjutpnZHhRjgVUrfb3wwZETFor36ObRBhi9Kk6SFuFZDrhGT1W1bxOmtxicTJEUtcPx+lo3
Y7LiEb677hR6lBM7b280ITO4uXlSdREIuSoKzPHyaXbM/oYglFO1V/ySG9/+zcBzsFkP97+lRCns
2mgf83yFceICdld/Ca4JEksOcee3Iaykw5O7yIWRUsRHmbUtkw7aQYn4qdc4fj1Dw3CkniAu23Xy
dEqllFYvOCgWEBGAdo7PBkRWWTmyDBzmBDg+dfl4cRHauCfW/2VHPMAdgHlkZCjyaEyMDPH9IuBl
ysBMA4tRkmrk03qxDD1ufHzHH0Y+/nh8I+70VMoh7XxdMOEyiWVm6ZNhOSvhw2GjJVaOmR+4krCv
W6V8D8b8Nha3476oLU2W4sv28jGKyLMp/khKKG26sMrn/9v1kplfeDlCj0S0pl7PuVSWXiE6f/ng
GO5wZMqviufQ3+zMBItTDFO+KcgwCi49CsxsixPZVcy0VCulGjzSBCQfOL0Z6T5zt2xrrFvHtqAu
i9X318quZUvooGneu8tLIdH6pG+LpGMQ4pO3SM1KVYwynvUPErcA84hUhD2FonAZ3LxPpXM1cvTb
GNLEtEdog/Z25UKHM2rOFcS3ybKdohtJzsrnsRPRKpwpAen/ex6JcXA7gms8qJA1VxbG8HOQX/3p
9CrUZyIzH2IqW8LtJ5OeU1H8xsc3NwQL72VItN/WqvOAmAOK7vq51H4FsX4JR7arMpotzPXy7o7z
z/hvGeQWnkIt1bcSwCM4Uzb+IyAuHO8Cm++cQ5QwZUak8d7/ZHVfJOvFA+cr7jKZzA1VSDis8LIN
F+z9q2+PWewahZlNUjnaqEsgPjJlc6J2oSzCimvubknj9sGMTkG8TN04ooS/bW9uSbdiiG/3DXoz
dtpo5qQ/WzdE+sgGB8qHNDHRO1546j12oFeoVehBw88YVtHXXpXrdxS42VzvfKotW2LOxhTZ+2YO
K3R4IXrEWuR5rh7JOzyX+gDOCXNalQCzkPJCN/n65sDvpQlQKYX1VMgmiYVUtWGZP+ncGQCryUjm
0tvmrNsfPxr7ACnUw50MAiXn+kPKa0LtWq6pXP3F6Bs2RF3vAljsPOUIKoGY+VMxhZ2bwf11NxYT
eT9YmklRw+b4oMKRZk+RrZdpy6bHVcSgwKV8xS/10o3slIGUeiX6wxrI/WmeCWpj50mC3OaV40H7
dYqLVz4etJ5Csy4wDrD/UZQJieklJG/Vp9gEnd2+C+b7PJRTveneYRBtHMUV7rsVodvAFG4ru1fk
3nncffaMtXUPaEkgU0IQxJ/O9x2HhlyHZnCUwOIwOhSNDsUC2gADmyqQjNhIBcf+znJbuZLM1PcN
Zcl3O/rpTMHkKdprGxYUoPRc+A+ZbBZ2xh5u/Ct9Uqh2cWAjvXnvWxreVglvYdM2H1OZEb05leGI
jlGr1ZNT/LxJShWoYj+5h6zYf/4/pd1QSdYFPME3jWMIkJPfSGpNCb4/S/PfrWOl4rH2bygAqJFY
Tixi4rMeZ4Y2mBpMg7Hsl4aQGhrjpp741cU15ZWOXVj8XaUSodlAWEs1tymRkMmLHCk4Z+JmJk7e
0EV49FIuQaw783Z1Quah4gXeauHRSggcItx1Jb2ZAdwmTA4DoCizGeZ6HvegncLx9mpD6Jkvvepy
+AvH7uBHUEiCpw4ClDmS0/8/QR3FM128PVlpF53LiZjAYfwzvVD5hgWM0yevHaD4i03E14hf+BBu
TDsDf43k744LjtrBuMN2sfZYKWwKHtbVGIomxSkxgrUBKwRJiqJNflhAPjuu48eF5akkd9xar8+L
vMUw0rOtplb6glpI9H8hdACjTD7hm0R9eIM+qpXkvW9iTLCl9K4tZJcPmeTrHOroOhjs5utxwK0j
O980aNC+ms2pvcOnxx4BDJhDGrT37Rl8XaLxeBrYdMYlXnzhvfv0agbmroGHGAUpu0cJtF5QJ6LU
simxqXIZdHHY92/RmDpAQmuRaGDGn2fcW64pohneqLn/CaFowhF2+XTHz8vA1lf5lTXqTVu6afdS
gCJHRPUqJyXqdXN/lQv9tGLMBuuXyz6PvCkUPwrEDIxLotE/D/ArtSX5F1qN2WGF9/+NWpWvh4+f
ApF3UO9hjWJ7ji11XPbdHy/GemjhA38UHa1uubHuBCqRDC0z9xmOqbd5vlX02ojipNfLdiy+y+93
vvm+z3DxAVvAjW6TwE3kfIzfMM+m2IeptdMLg4TJcmaCfdxZ+4+G/TSaHnvofGfjsmbSAmUaZMJa
sfK9umEarZBIyCU+hrUPeeE2IBEZQAz/G1MDalmFYZ28KFHITz6vjpvv6tQf4RsS1aFp6twgxwDy
xyCfcTB1HkIe9eBXHrg8GF3+OzSz33sxeUejwErLiGN7WO7uaexmRWGLmMsH8JPx/OTI3MCnOP6I
xmdadImmXORhjYHYs/nb8RWEpNLIyK7fgQ8xo9YA8ag5T6c/tGrDixic4UdvDILcZJCD3EWdN8cd
HvDjMHYarf+25PzMaLMVZl6Xs9knWQxwWCvRrAuZHxQczdI5ur06QNcauE9t6XvPTPmzo27rKPLk
rA/CbO9kmKWvWSw8MtiGfymVuZ62uUsE1isYbu+TFFJKqDoQ8ecgoE+LjwOO3sevatrkGJgO+buC
5ILhzW262+hHpjItmT7XsQhJ5P9O4Y6GIvZPw/fT8lW3SoQz4dZQ2YdhK0rvHDiI40ApZwdbxb34
0zVt3UeOPZsEEXr+nnmTm4gcBtZDxJag2tPe7njqyOfLqxjB0H0YRTNrFutnV8yF96/fN7S09JiT
36iTxBZHQChM4+6qOgb2zYXDq1HL1Fa5bZv8igSctotYuVmsq/aGTwvV9ouvW0Or6CWZQd7aXmHs
to54A/hAWLwGRepWsVUt30a5P2z/e1PJ89xFuwrqgr74aM3aCosOg8HmY3QvXd9gNtm9XN4Uuo8O
Hp+XyjqoXIZpZYwJcKaklD0C0UihCFCWd555BELCxPl6Zc23bke2VmdWNSKO/m8zwr9BF1rHDj9x
zrbFHsk9hwCmK2GyonxP2frcXEmYc4p+hMpytD69K8bB0KryvqOf1Kc6oy6Jm680ZnRrqmju4bz/
JqLfla402fbeGYQqGy1cveJ5VNpQ6M2UBpuSI4cdV7qGVpYpxvbaGwWxJl8eZWY+4Ygu/1VU0qKH
iyFTABE2xFWd/9EhKLe341E1JkVRZMMQaT+KSQYDW2gEsOM0k2QlGxNKd9/+l1bvJydBlHNW4tUu
3iwo20IvrjrvSPkDeWbylf5bclK2e19lWxGgbbEHmXqkAwTW/yNN4pUvcfDBfcU8+snu6op+/fVP
BjaBe4nEbk58ALV94gsrnKfsmzpDirGZx+s4h5UaLOQ56P8T87nLfjXtAtsDYKhNgek+EkC05yMt
fTltNlTsqhHBdVI/aGmTZMSQXA8mUjki1nQZhfW4hcTHzG1WhL398yDQHRLfVk1c1oLlcyQiWD75
HVvtKGSaoWjtY2lo6Idfp+GXd3mcn3kmSqJ0gGbXtV9g6TnYZDZi3G/dmTUPkWsqDGK61f/mTD5E
tkNHD5J3e5uNvPzrK39OLJXdO0nW4ANd6quAXcnzpEuyZsG1E7aE+QTnCLCYlpnDY2GjtNjLCN1/
yz75DoGSF9O/4IHtmbdoh+hKK+Gt9U3Frmnc8ZRf/vNvYsvaHG+wnaZtIrXfKrkEPTz8wtd64ldM
KESVGvjzcueflLkAGhsyaeeyuAZCfvqH/VYIDS7BWRWuY+dTMjMH3c3y62ld4Q6Fk+czSOeKH4Pg
ygZSul/G6p8gaW+nkrO5WA7C/YNIjVF1Tm7mDTF7O27F4wBpgtLBEHJveT9imKffJR/ZnySCl0tU
lKKPinlwIJcviFMmaxlMZ7hXZAE5qe+crB1bcEwdXqWhyJtUSr0n74CcK3XO62L+OsHF87YKwjIE
zp5UzqJmli1bUhsZxU+Uv1rSQRbyNX0/kTN9LXoJjjAwEIQdByu0T9ieIRfitGsgEXLLm9vhSu85
wBY+BXWkh0rTOZkEgMFBdcaWerEUOlc7/6VLxVt2Xm6lktaZ5KLilhU/IJQO37FmZg1XmYxlx/4E
6xOHmSXVrqVpCou5RLxKKSa2Nw8p4WIJ5zY4yYTAmYZCWnQGNe7NXFq5mfi45oZK9M5zsVUvVec9
rSrhXcOnk0pwgT2c2SHIT+pJpj6W0WNfJjWL6nLARj6rNVFjvhVTCtZVg1RJKUycm2q9Dz5qBiHd
DYheiUg4C9ktLwPl9rscbTgLn3Ap3GN6qgL+MTNmOnE5GoBvPo+dz0Qs35/VVt46E5cH0Vzf263i
KYh5gE6FHOxArCiTcDZzJ72Z7Ug6GWCPag14N1vjHVohsPxxu8dT5vh5gUwUI660J8M6WhkRAX8N
ZagYXtbz06N1zrtmv8onE45iIvR9kczR62JhoH/hjbElCJZIkiL8QW3+4gkGeOV/B/W8IZ4xWQpt
FmGI1PCvqQ/d5qTCueJgHgNxjIQBAFHfjyIi37T9DNA52cl5GrW0jmROBXn3Rh0vmwnG96bZ4Wo/
Yn7rpEZJhOakSpdeveLWeh/Tg2ZQrTTfJa4VT45OWciNKwS2rFGF4YbMu3rjlelwCpUEsm1OzkbQ
mQWVVpByVZMErKjTpyKbKmiMJnk3kM09FKFn/k2PT9T/Ohfjf66D5yfnl+DlzFtGTiPbosiKE5Op
fAqBeLwJziW+fTrRCwDzot4afOkBTOSl5EiGJIOHLE5jNPobqlc2AmNqodzE31ln+a5V0JoWPDzo
8GBoAd/V0S89JtqatdEchHbaKUr5vT615Z4OOt5U59eUYbGoEUpo4G9yeu0WSS1ah3kQmKQm9oPr
NkYnua0UbXo86bTWq12VbIcOE6adbf6vVy3Am8pUdPQkWYXBzZvcNU0RHFmz2xEG2GmwK6N10k5k
CmR94w2tYNqbivkSQZf4IrtbIFInMEOgysFTTFRO+KDP9RbAemdyeKKeMwiajHEjUVPX3hl/TGtf
x8iVZG/7iUGf3V4tvZVbW5N/MX63HqXbyd8YzS0d07iPypjN3D6s99YnRE9EFYctEND2vFkd5qe1
JAE5jUP4MDBvb6GMH9gg2xzOEjsUdL40xqu9Z/Nv9L9ET+AlGmZO2dmFEzadieJkavrcb3bKq8uq
WqnQc1/fdEs5xRexSZKiFVI/NzEofNFrIcc6MW0a7gWqCm4Jaq2gW4tUGeBZfq3MxPa5BUDlFW8s
0+JRsD+Ru2frT8M7ZiRnt6mWX8a9zuzHWprnKyOCscvio0AsrHCmWoPKL/qSb6kDxVmLsMap6VrQ
IQ8spYc9q3JEDczValJqt9xv/QljtYC6RiE635scO34Rhj7k+LPQBhQt+ni4vahxJxFHjb7ZCUBE
rv/d4/Y5WiJQ0WMgwB/w/7IpeBdOXFlaLNveFlWi9btiDConQWde5CSGOwke/Z4dkveZppfWv8Gt
0n6Lb22dHYV/PLSB0iTdj1EnpQygYlRxjKrTjF/81rE4aEVA4B/sU0Z72nkzM8AoScpZ3eeOEeBz
aGzcZCZ4gwMCMC8XJs/gtVgMYVlK77vFVa9H82WOMMLHCID8EeCy+suZp7ak2mXw10eF1JlJMAz+
eVFT3wJ+ci4CYUjy1+L+L4QvBGflbyBcIJ+4oZvnUc70XrKiSxRChtLuyUJdr/Cyx6Bc65zOpNQw
538cQsxnEfaWX9OP0+CXMc/alpX/kzHq6rbUlfFli12G2WyCLPltup63+ZU6wdu2Xvaj7l2GC4aI
WrtUM+C77Z03JVYilRrHhwN2WcM50imR4d8j7Hd6E7l84IBFNrKe9zOg8Qk4/4vSehGLolTOztKX
Mlb8anzIupc0M0gQCHf2BBA9O4leo1gxKj9W1zeJxaqLRpMx+txLbDq2Vzg/KR3Tn2ZhICKbFs9n
tjBTc6AxdY5bdV4OTtkc5bsxKzhZsiERhz1iA5sHPsC0AbLHeTjV3HZH746xe1jlw6Xp0kFP9lMK
eUFvNsEZtJ8jNBrwYvQyPC3NgMoE7aIfLYJSa42XOA2Kv4Kda49JfmoFaOilO5lJQS+FWtkhP2BJ
7tX13hruVXqzdmOZVh31DMeBI+yyScK0QCcMcg27vxrVHisWvNiGvo+KX9kWuvUlp6fySbgU5IvD
qxl0F3LbzIDY7osahr9uJxQX5HfnS67xxAqDDAnMQkLxCj2Uzprxtgvf2BqCpx9svOYNlNNbHAzn
8y5I3MTI+BnjKWr8Yb9wr2vKtdl+E2BguM412N10weOA0eWfsCH2WJ/0kZoWUSmyR2cQaiHMsIJ+
0a4YB02cP2cflhAGKCPDFQznUUaqf9+rI/olhHQAMtTxsCU+0eGno/kYGcOXhY2MWeayUk3Y/6+w
iwjUL0eNZXgGKD+12q589omqLRZ3P1jVgZgF7oBWCGF/i1XLTiYB+lOSB47DtbbAQdftlCZlRZOh
J09lZ9Q5zPdA46/kfb+569+9p/f3aaZ38AkbjkW4CTsEzfJZY/F8gS2s/PMxqi92rxTSkCtF4wFi
PBYz9407mYK12bqA9IyDkk1VVx8hWhkLChur+zxmkRUKWpvC1yR8IrYiSJ1bJ6ckQwpenUIx/lRD
gVQ5XZ239tS5gjTH0jA4tNaI+KYjFBrpoDnX5JePulSebLMC7l8WcgQY5Lv2vwhT8nH6EVMmzrHW
N6SZ3Nm/xYSug6VP3+5ytLwZP0gjQtZT+6+++H9fAiM1F/h1bm+jHmnLaY6wDxUbXi2pHAXtIjg0
ilAAjZXWQjAtFthtix6ggTHKtxS8gFMqRebehadlJvc5LxznYtxxH/3siv7o1WXF77J9/JPPdwf7
CnviubbYT65JlaUMPUaMd7dsOdNEiOu55briiMDZP7voKsD7jMMFOH4AO0N6WW2/2QbJmYdZ2bz7
CxWgZPNllFRnuRMpAcIWv3tQn1Q1D9aeEqJMd/x/V+pk8WGg1/kXIiXoOuFd27WqtbKZxQaQVvWG
ma5TNV6oj+c0IjXzDgQja74HT5XvRhXrhO6yaMe1ByhTj5oY75CVDSw+iVYasLH//k3yS9jiLCbJ
w3EiTnuYUypP92vT8gOJ3lkZMdYBejYGDkbIDLGvz2Ka6e1P+4AXtUBFiDSRb6LsNR6nzm7sVXwo
ptOfBp2NjuoJKe4bc68K4b/o3C6wQD1m45xy4XY7P0KdIy+8t27HXYcxCeqJ73oD2hLm/HtFFMfp
emwvSv9BN7BCoZpWmz6jAZ4EsXSDRP/SCKICOJBW5/iKwBnta4oEFg4u9cfNpS2J5QqbDU5UUid1
mhEJw2kqA6/AzQTli+ciaRJKAs04xHKFq4S07gUOsXFg9ixBMpHKFs1WFzajqAm8fvaC3qZLpZLc
k5Yzl38O7JkukoimkRrbEBk6ds+5Oa1ccFkEzWRHZhy50A1KEu9CJWVedrf6/7pN2Yte3l+/sOQL
ocghImME1NxwZ624nRzJBgBA5DGpKRYFSO4Lpu608dY0VLgexOeWY3TJKpDziNGxX6+HP0KI/zTw
Zjldzsgp8+/Xq3c6OqXF7kALdwxZj6juQKgvJu64GjU/3xldDW/CQ0bLBHexC+wtyc9RLgiy/YJq
rUzctC2hE18Ufl7jzTEvjbAJSR8FfQcUhRMn/N4/g2oAhAKAMgOPzFIEGIaLKMxBmSb6CScCxj65
OtfImXX975bdvnOGsarSMNu6AKg3YIIiw7J+tNjSN+tErA3rFPg/2wh0A7WKtR8JWjWBOii+SlWe
UYAj/3pBS9scNvVWWXqSkjaDdMDYOx/H2mSCsnsl6SKpyj2Rf8Wmf5864/227e2mK9SC7x5mrZwM
Bf/2Kr5RKm+ov6CoiSuxOeU/shKwOwXPNeXS8rGGV7xQyAEknMu+kt7N94dqXay39+hAmAuZOy+0
HzgofBXtFBfAr+BASmlAD/IWRiDAEtG6Vp0hOl4YKNR9CRaouGDD/i8Spb9y6IrPuMEoW6BQyzJz
PTKi17vHdvNfAMGYSHK5fslGuOuiFgUG2Lvg31KK7zXA6LdaBmBFbciC5A3D4KSH5MN0TPr9vpSo
Dy2mkOBc3/p5Vls0LFUb1aE7BywvVw0lXEf7FBj8842Abzj+5sn4WCGm/uAIq6s9k5nG7agTVt0J
83ANPb4xXUY17AXFp3wB6HYif24tWQYeSL3wc5KBzqRARxpAOoUTt/wGui1Dgr00RAOEbmfBnhWT
pFrOaWRPyz+8mZLbLKiI019MAAdJU8oMo53zFbBwLGSQO0hLb0n1/4JrjvVlvVrBof8UDxdgeT4q
Vc0ca/uNN+6y714HUATR+P6+raxgmPtypfyD6ietWyJXVunfbgDAnBNQAza9WJf5PRMWSQGhH8ow
4U+/rHcZFG5UFWE6W/+2HdhFKQCc46BVCQQor7jdHtOoSP6xWAwrPuKy1Fjg9Ka8O0VjUtMYszsn
zuzmilTIreNerXI86R0n22YrRuzCLuOnGTnXv0n7OsbywSxBAA08T27L/QTL547n0Crbngy2J85q
9HmKSLTf2g9DkUPSxoQGZGjKleDWpTKGEglupq7nIuYVdMXmRj+r69dhCOaKMgSi4tbo/Vixdnm1
PC6iK2lgURrvdEuvEiY9g7q5sWEAlxPT9k6CdMop+4RGRWO2QYKfUVc8XwpC1qnimYfp4Qd9RFPI
ZKtlwvUeiBwqXRsfM5PzLROWLQKXjQkvg6z65UQGi6LY5Gxe7rbiPs8IlqR5VFJVbi4HPs4Ol7qX
zITpDRxucUby5XcfeoqrZMwwTSbTbfofVj962nwzpC3/gIz9xKiRB3ARqri5GRhSjTVD6xfH12jQ
zs6vXhRW9/DwzX0bNfXu9ZZrVnB0yeWUEWKGWler/Wmr0iA1omdDV1EhsmI5k0zf4WWIUsavl4dd
zczy+DCppB2DPV9I77Eu1bi05mCjmwDstr9si6NuD7M2iaiK4VliKiQdppYbbwUrjXOcL88D0gC1
9tyylQW5Jon94NbP5ZSvRvnW/sSx+9eycg+R+UEc/k46YJcTbvhx0vfcpMQKV8pi4oRpa0TubZ9F
vQHQA5SbghbmL6TfLnS97FTRlM7EMJ9zqY7Dg3hzo9rxd9C8BsDH+bi0dda1bPXjL19CSICMWFDs
bVRbZa3YMPmP9O4yB6K+np9nKxzOsksh0gk4n4lYl25FO1MIA/WMgfcMbLBy1oXVizGxMI/S5TrI
mnTJOcNgBAYoUFDntVwAg2YUaBIdhpf8S9NufxVMrTBJA/p3rG5v0PlPUcP5K+/hpTWQ1TwenWDy
ugyvj/Gt1KjtM/BQgyCLiMn4g4g/FBkw+C33YXmG+qYS5sJzXooSQRNsAgbxnKLEbh5R7hqgooI2
zvxZOZDjvKN6PJah9kuz2sDLAEwASjWp/NUgMJko8OPddvVRvWwgkVsaKtdOSG5A6Cm/L0he2JT3
v6jIqUEYeMdMc5dzzQl8jiOdJq923PKn5zmt4+hwtkbKcZYb3V0jVcEHMSMeNn1yek1WgNGd0yTD
6LTuRneGu/tfcqMrj9KQb9eY/9M1x9cMi94Xr4OBhsnbyJNviZHOtBEd9HcfnNgYx+oTrgUN7WpT
/CTDcj719ssyVixvBfcypy9j0rPswQaHhiOBoYutUs0l3xqU8wMOzcykFz7HgVEEZVgJWzFhiCgb
4PnnyG7t9JbbwKtqsNztydIFawNH9u91tNDz0ygzpcGlcGGwj7ZTO8REok0oDBEnsjwV61jNQtRR
1DXPSQWmo1EmgE3ikToAAGdkJiLHBUopgFN6wjzSHf+c7THF0z9U9beApkX0oh6dhlm276OEx2Th
e41GxPakypDzz3YupDGge5czSxwyum+zNevxmX3yk//4VDkze0bpzPQLUzco1rAXr7kQiukSGlWm
aiP5XcgkcG/mM35hjLvlakgbm7BZBHMf1khwDpWbntVtyy7+3PUlS49uIFfZNM5vZeWZ/d6vj6sh
k25/+n+Nu8GzOFJ0UCDSnwr8Ne8NoFiSyluAK7CLzc/+URA41DrdjM9vSDozPqBZmNc7oTC947Ha
cjSxSTdiMFeio8ZwaDi6/IAVSXmBM2DoxPgZC/zUulzt4FLWUsX6hjBzq+Trs3++J4o+bLSugGbV
K/nRYcTghIpSb/8vcc5zHF4PBNRoau810ZLJIOEHTTitnL2IzeT0Dlf78VlwiM7BKyy9iVb1SIQP
c8ViqG/DVHiZuDvBpPT3e6vaDV1BxVutQJ95EawaXJ6PB8/yhS6l0o32+iByGWpgOpgCsrglEt9t
O92Zp6F2iF9Ocaddz1waW6DnTmJPtvQdBuu0XtKDvSNvrglaoYi7MFlAVzxpmRorYkV3hesieG+/
jiZV7rroxa+ai3sJTCQRIilaUvXxoaaIyQWoIpEYlHnmmIWLL3VduhUB0eAdVNQbqTjym/LhmrOW
Kd3+u2KlnHQy7tlh4bCDAnbwjOQ+dw01BdlV14L9D3MJOqJPptHwivUoHPcEOCO27hZslQ7o3wOB
zB6cLGQv2xObi1CnajoIip7ddVhgR+kPzcKOiyx6e8QFA4C/OyGghrsz961gUwD0enZn+MmVAP9f
+i4KgGDfIFV17bcObl1kG35hmn4ZbzF8kTsTc2arkWkQcWRLJuLjABzU28B4EXmbGweCSJVl1Kyw
qw/TBDm00Y/8nTcRg7OZNEXoUMZ+2QW/prVX+COL13n+L0YiVsbxU3f+SVhmhC8Op6JQNVFsVSDG
Du9AQyLFFqfqaa7NOLmP7gfxZblADeuOiuvw5Qm5wsAcRpIeMLQIE5n7k3vGrD52D6tv4VPD0LEk
5VNuyi7dmEBKgNh2B/dtxeUimBbEMppLuDqMZFedBsg/Vkapt5UqIE6R8KVwZWwZ6WzQF6T5wyFy
M5EcRsVGFqEin0AkWi7QyPCd12ScTSZt7wJAKtOAYmZ0Bh9kZVTN2Rd+ssu8rWI6iEIbUhzKTFxp
pSTxTj9kE3p226PfYOwys1U3iPsMgCsCuMPcvOwWN6s8eSPZD8q1leeLyn7mCokGkeT/bTs7Enzw
dZlI/ZQ6dAWhm23KuKzT45ocNF7MXQ21LV6mKzjIZwe4yxHXnvA2bPjHVdL0YWaCqZ6cyWSv7O93
vWiqQ8Elbj1ULlI5bgZpsDt5UOFNhjvbul5Y+qboEc443D4VrMgmjYPD0iWkq5NogaspCWqZadar
A9RlqQfC2JHH63kIQoxwOjZ2WQnz+biBNWu3qOpb2M4VEWD8wafwQKKVY4TIBVuww0m2O2Jcv6hD
qg+IkLki/1w4+dEHhkh2lFy4DbivX/dBpj7omN/o83Ayyyf0uDDl2N6AVZws+c68jOmrnu9mhAOG
yhqIGgen3KnEc21RSx4kli/hO02hg/rJwa9hEowEm5rcapD99OdoEJhYEoiXzbGtR3jX5hYZEFTq
GQn0xKFD0GaUk3dla/45xX7OoBnqYXVvcL5gwGjIhwcF/ITSg3Brk6H/Gafq+AiYjE+6ne4DJL6D
5wBDqWotkJ1FFBvJ0xkmteHRbccV000ce2MUzsMKca8k0Pa18gWu9Xazl2MezxAryhaW0Xbbn6XT
t6H41bLoU8VuiL69BceqTm1gkKdl8aEt/hT1/e5or3rAW5HJ3PrYWks69ngp0fI6wC5tHYO4qlYL
3HOmG25gikaexPMuHxbt/WXx8MWOr5gt9f2jULpLubtILNr1MNr0I1jTsFJB23qHFV32l4e1ZZP3
GqAbxgZet2K8N0bwF4f/rNHUYnMNas3lEhwpoOXMn86lr3XHLb0XYxNhtPX1Sl6ohbVcIdpFf+33
smzJK3bZoWyMsnuOrJuAFGC74vDHDHlzlZSkOemQY3a504KSjlyxq51KlzVimqBbqrQFZcwpa/eF
dXL8F6B81C9K0gQy/DSH2JcSEzQ0zqjSh+oZtdKersrZ+adJQDP12COWQq9bjZga66Xt04OIUWMb
AokyezjVIewBinMPxS8ZuUl3jzqwRYvxJn2eD0gn/+mXEiONjm7e3eLuh73yPuag5rkoVocBYKvR
Yn3NqSCf8wTsaBjEOfm1kfGstAKEx8G6w8EOIxbg0QIlliq9ElVIK+40N+lR7g4cMc5Q1+NvxSVP
fZr8XxABxA9JSuBW0QgIi9+LhkGUL44JzBuknjU8aPHqvhTR1nXPkIIWXAW8D7oGeXH5c6ZeQ5GJ
uxWFxM3ZoyRBaR1xaY6/mK9IA5fiQ0gNrsrkCLuxJFYzFzROIR1lGNrONpOiYyvMKjvLSQlgaozT
PNr5zMKA8l2wjpRkJGu/7drNXKoqKLwK26pzXGmvX0MEvhvy3JooFdNMiN+rb8xy18H4eKD/NP3M
d70S1M5S8EN4FmMekCeB8apnuADqJrFE1DavcDDMBkg9wdUZ7HJcSm1yIEkXiud4/psBr4Q/Oc7z
ZUOMNuvKOUb9SrXXOrYYYZLw7nXGDvUxF9UP1wHBvk0q4/DdHXbg7IuYDNctk6JyWye+ralozwWn
3HX3UQGA75wt5L0IkMkSgwbHuviUZsgyjyJrrvdq3Vj8ySJuv6Bz3Eavs2XsjYY01yyvue2uXlHi
JRqWhmgg1pSY/cXGMT3diUuHcmQlGHajW+sJOt1TwG4vRj23iVqj/+e5I2Su5Iv11SvxUm31fl21
XSXlcPjuKcF4duMVcVQBo4652xi39kEOGi625RgFRK4QWXPTMaXmEnkP7aqg0cnl2Y0t0Ius08r2
ilxFLHmsDCh2RYhtH6QYVhjI2tb5cWi1Vu3HJqsl8PQaga1FfEulSBxxbQNYjx0G6WcPXw5QTJpR
fdZw8vI1ofmJ/12Mr0UVICV6cyP5E2u6wqe8s0PQ7QOXzAXNFUXtLzzL5h2Uum8oDWrgDUBMlfsJ
cyyGimdLNPbwpStaT7KYv1d2dvj0mpmZfq1DhSVP2kJxAdhpDXldYzE+PK7bZDMubB3yI+TzcMA0
piUcX77e5zYTF24bycOHsazTb422NdqyqSMYOnGtz3INh0qgZbSxviW6CGV7KBVIQktuH+f7Hf2X
hlSh11+Y3t4bg+z69TQmbyqg3y/3Rf3q2ecA3xjcFdiBx5b8x9fUees/DOZ8vzlri+t1ZlOG1T9X
I1y7OujeCUBLLu1s45BASG5/9tcAJPG8NAooOVjW96+iyoG7VtXJn3vxKEMK1xD2DWbkreZyGJ5e
oj723q9dz0/T2R0zFFnn8QJIO3CrZcCCLoAfJjmsZznDlJaNJnjtBUVHPLYXmIIWTK9enSaupu4N
uT5yeuq4rPFIjrmFzwGX3VT03V+gAmTSlbmPXiWFK4xeQnuRPG6mHG2UM1edZojNiMbpsXfXHJ3v
YKuxIic6S9orA8IecjZdd+FcguL6uEukOMHVdQifCS0eLscC3sIwFQ2X/4ysmjwudj/lvd6O/f2t
wXPbTKveGy4Z+vF0BuOFvCcAxdETLyiXHGhs1McOQUSyPmKomiFr+IS5WZz/siL+hLsuWam2qouS
CeumAoeiXCn84M4Ylh8g2slHdO0WbYt/mmWGhA4My2AB72UtdfQf0Sf2FKvsAqt+OxSGP/AjShoM
v9hVF4xMAAr005+NO+PVStDs1k1l3acQPtbqhMICuwNKSjBRJGiiobSaOlx4Jo3MIZBtRPuiR9eI
skDuJE4F4lgBIV7jPILnVbEhmHxmKYtiqSc4NvfWJTb98LX/dwNzQyT23mWBzsNmDi2XMc5hMoqD
FAQeJcqX5ck1xXd15ptAg81SdHXGqZZsjvPAjaMM3xdl7na2TLXK/U9jmkUngnXc8PbvQ4ea1kc/
SPGAxdyAuSa1BjSjMPmFHtrDpg3BPQT5+otforYvZAGlMJ/JM6UzsR8wTKHEVyZQjxiR/yFVlaWP
DSJs0T6ySsqAeLoxAWlZYUYXYRJmelVl1wryZjZO0RjEnvv0nlI2kyC5Jn3ZHr0cLGui+swIumDq
GkewcAAA7HxtX1Oo8m+JzanhsinAt/dq/uVQioIZ7HMgwPAkbnYyEzeBcMdRh2O8Rfce3K/IC39S
KqqxU0fMVAZn0u7gFpDzaPf5pwkjaVqdxvN7z9tgvMBUHftp7Gd8VFqaHf37Bctl6mPd4yl2pCzs
NG3RwI9G87Kq98cx6YWMiOvAxc7lIR8cPQZ3+GM2Zh9jL2tyP0TwVUEvBqYhHArpg2QkxMAvZtZz
ERA1ozu1MrZ/fJ5MiyfM+AlTosjVViHaTNpb8LyHUzuw8IJWdjGReBXDbst7CBuTEbKazvOLutBd
1+i58owW80rrPhNrMTWPL+dBIki6gxRkE6qVg9ZweKh2T5nxNydGKz6zW6TC/Kj6nsbNrbE3xckb
PPKIZ/kJ2rBfCvkqTcIKSoKVom0lVPO7Fnp1Cgir+j7jeSupHSoVLCEdu9RoVZleYxsJtxs43EmU
tCtAD1zyn/yH1H/q+sO7rqT9bvloWfqCwL9OgBUsLoEI/DDHUWcDy/s4ltlaFNp70zD0GjR6waLs
ryadCjSKCoezYkQbHpVov2l3fXFyinwnP7lOecXYGBPURrGEdrVogYIpjP+Nh+46flrHo0/YjMxW
1tGxH+CW4lp7U5eFk7MLhPkQxa7cnKsquwNOOM0uIbv1pT9RkAZqdqY+yZXIh89H5PTbhEF/WV4H
CnhI4HznOfszrMldk5P/L1jzpvK3iNy3b7oLREM/VHB0zsAsYivRXRP4Ti9gD63lXoNw+MvnLIdb
PY16moGztBX9DJP0oiIE+zsd/uHuoWFJSYDLRLWSn1/f8Fiy00MapBnhuGD7lSFbs1HOdQbS8Q9X
6BkH978qvAslleuVUt7eVmpSWzKTP/9ygZaH7Qn0OQgONg8AApzH6EOsHs4FLjJwkUjnOMp5ZN/5
8K2ovDWmKNj0vQyrCo10dncHjIdLkjX/clLvm0WG8dSqIZTiw+9rVVQFIoXtrhanphZ45Fygm4mb
fjY5W3J1y6gagiudRIgzHGxKYeJRYcuL1eS60j+23uO3OAcy5A/CB57Kv2Lz8si2kVW9gKkcouVj
ynbH9uadnv54bINCVEQ9vkXHV9YuNatNhH8vwu6D0VoY48D4qZuj/5yJrbFWeV/zYy5icbdhznxB
DTErGDFcFmVeOVET4ScqIevpY4RiMEvjHLBa07vniq+vXhkOEjV79ppZkQNlheDqUHe8QDwq9jwo
x+NubVFwCZjiqBkiJoOeSv26qxoAp3cMoxVFDDDfP0PPrlSdr4WEGC6SwBf8XeSmhryav/kOD3FI
TblAOifsrIQlEi2p7AK/q3UigWpuD7KzuXSr++hWp4j6aiRo0UuTapEEIevA6ru6+f0d4ojkyLG9
Ze2hIU1h8aCaa4d1VHGOO1oVpIpAK+BnkRFh+nAGevHrTkpXYl7itpl9A517dNwIY3fXcEheVR9h
LezCTkVksCkRU8cvRM41AoI5lNAqau3Ski9qdz+rZTZUBOdc++J/7E+YF62MoFNuUXpeb/P2Iv0E
VRXw1gTTVX/6Duv2Ys5PEFmi5MX9+4Ca3AMtUlWws0lU4+bolD63cxwVr9Du8OwPFgqRDnktvgXA
4ASxI4IJAnTmhB9Se9WfUZXM2f6EPq4NSWDEFqoIJmHX1cAT8Q5Dg2GIXCWBCqlFSmjFVmCPjIRX
Ll7Fe8wrrm9m39V+37HN7L9BLosNlIfEO084hCA1OEnVbnFbpd4dV7ZDC4C0VgQXa1Mx9lcMzDm+
isobfiB6XkC33rQ6T+r0fL2f33Y6zYI0TEqP8Z3HjAArH7f67oadBUT3gc0nGTxNZeOMPzbOkYxY
T7k+PO60kXX39v3XCyKxWknp+sVNDQ7cQpPG0YuWcru3lK+TrKPXdGa7p2ISzTsfgL2puyDN5skC
aC+lsvEtruz1AKV7G0c0ZPYnrgACbq5XPIEsLXECUCqyKn9rFznO4N+V9H6QDgdHb0DXZqQN+lzc
7WwWAFD75ypLEQP/ZZx1WSmuUes8Cq5en6hp1bHMBRHlS3qsVXyg462ftrxG1KI0MqaWFEah4bn+
zvh0rhF+wk+Vwb0+GsSlmRKj3wGpEdrGRYCdotvr70zoQNRFKuNRJlyURqajaqDsZWXzfRvN58Do
CmqnXJySPGm7KaMNNIxcPjzr5nJ93v4wpSMuXzQFsrldsT99mZcrJdJOfDNvcMni5EOk21i8ilB6
Idund5DtONtfNHoH0pCtbCChd6bRSLkxOr1J1XsZ8qJgzv+vPH5xryxse/x5QdUyGkKU9MrsD5qt
J4LJfuMKdTzxosjtx5K+TgaP4Lfqol0YsPN7KEnLPzo5gGZ/5jW6MvK6stzjR1EXuvdIqQCAguqB
TSTN6Y+lEI2sR0qlAtXA5xLOpy70UjEkTLK8a1uy2vShMHT8NQbyEH4Yos8noUxTswPp1oQrwcNj
P2FSiD9MPwnk5TrzsMRilZCsBipW3jY3s0b25lZKli441jT8n9nA6jRcxEx7w5I4JTN2ecPEJfXB
+wNRNq+MU8JgRe+1ygE0h566Ir0dUOXOwBJWUlsiWAWNll8LvaIzd6VaSq9jvJooqBStOaogGyFx
XGVWRvKAI/d5KBgXMVg+MKsUSqOrEX3xEfRbbsIILFLb4V7zKh4wSJDHiv+a81f8hmARftlsQ8Xg
YA4ymtrDHWlnkUtlB3k4fWHczLY9GzrPCkyrW7VGSipAHIORJ6TOV7Dsrg1HwbrFOKkp3HBU0O7Z
HbDERGh8Qz5NdtC3wbQ4n3w15dNZH5pKSBobwfJeljk9wyZfcRCt70e8z6C+CePDtSKNR/mN6mBu
7uxyYHNmuTfR8IRpoFgtfeM/6jIolgAvLyXG9YymsL23InjIypca/vXSaY9kKBlNc3WXzI4TeM9G
Wivx0YOxu/w9kYgwfxlON2m/LFlkz9X/Xc29+9KpXpG3suD2L3meIsJFV5V6wOzT6cUmOlfVPHor
Z25Sg5BIw3X2aLT/lz7hhJ4HaEJpNYh8MNcfKHHG2KCGg5b5hi61Pw8B3Nk7P/EvF46/AFjs033n
voZKbIEmhZ6nO+ktUYEA7mPejzByjrJ1eURyBMbxOBzTcQt+Hx4qTPSk4kn86MSmiL85AGt+8Q9j
RsWfbeYn/31J56h1QLHKqe7w40hn4GFfYMYT37MRAKxf3T9jKbgUGzxS5J7DDJ4u/oAxT1k9cgpA
A8VRnXnvOIM+zM3pSfnNu7YZt5qG59IC1tblz2Z/R2eDl/DmXA2kQcnrMigUjyLAwRdkNixoVtxQ
qYtfBX3sc5BFQvll15QpNwG0mBCJ8W1dsTagKpWM2mJ8NmIY885FEXQnTACf565Q/5AVxHCkcpbH
qPfxwyGRnRfXnB1PaoGg0mHgOm380We8brItfiH98wfDyHGh26UFjUfX5gZtNXntV40FAIi5gt76
K048oLZM0BYvttiIdyq6Z9yyo8kI3IhfZR1QZegBL2VnTtpj1tFYhs/BoYJ1PusrPZQmZ1QprdeU
VtYCD8Aoi2FCczk5fHcP7izCUuNu54rRd7COQvxIdKBv0pyY/T7pt8DJEerXluyaGQecb6RozvBt
Me76qvk8mKzpi7fZikWR57Z0JmEUPd3jjuDFzCCEFXP7CuKApW1YxnPO9IKKBgTQGMTcWNLn5IUI
EGCCQ3lTkg6I2LUmAKa2FRWcwUL7OA5XhLzjWA7ETqKxiyuZHdeEPPiLdmSEsN4KzSz/6pV9VLFC
qGKPuggZh/xPfVSSFeKDSzQZF6CqBQB2Qsh/J7zdmaiksDV933wohlWRAQbb9Cjf0YB2U9CzgCqp
ah9ceT6nn2iw1XoSU9d2ML1FrBM2ZN+5cCvUnSU0NlvhO0LJcx+hvdZJcBdbwocO6PZ2P6vAUxzE
bOaX1Ka8nfFRc+YY/J41ucDRSMf+CBpvXN0ZDvyX6PPpzj67f5IeyXx+86+GQNyQkc4AIBzfikbb
RuaHsVbjcK1Un8mOJPmstFd/eBtpwe/OS5YaAxHaLJ0jHi7hMvEMsCrr0Y3EJhuDRX5ArCa1ExDs
pFKwWxBqGVnTHbXOS0Z4EIL1FDbL+bJxG5/DKRIEorhx0PsXRWpvDx6SUuTok96evrWCvd+X1h4t
DgQOzEzzVoFSoqgX9A86zd65HB9tU/h4ieB5u33jPBAHvpshkUWujRN5uGix+UANKv8LDcP5wQqo
S5jZBPCdnSRvRmXbFN4f3ogsmttv5gtQg65SmS4R9gJ8vnqVi2xJkk2zH9C9S7Wi+9YktwdW4gbB
tTHUjk5i9cOfvv7SPrUKUfOe5+NY6yKdqJvdjG1MwbgAoCHuf7NvWcOHeCgjRpxlpJcNm6jRQnAM
67eCe/gpHQUKM8fDTgxSrGcZ1+/ZMMPnMK0SUtCmQtNbWD9LekuLzgTGBKvkx4iAhf1SWAdiWRbk
rwO9as/DnSmB6tEl0aOXGVC2tJvVMikLuNOdM/wTUTuDi+U5EVCNBr28oT0A26Bfm1/v8Vg079Lv
gmIC0GsRwiDUpDRFr28Wz6cDctH8p7J9ibu34MIRTYExvUBZNqOtLp0WMdZmZse6CHGoTw9qUdES
tOpDpYgzPY0azzUlbHB4EXckO2mv3Qwn+L52i2azbetNGUtdFziDVV5dDulh6Ur66ZotJlUSvqtu
tSy5/+1LFtIpkSsgZmPiSQoWRXxJp75ynV/2lMwRQEuy0bQ5lz6hQtO6hy6GHRSfVpZceJ0HOrIG
jbL5Dj+xp4ngaZjOXC6A4i/1e3H5zKYZ/3h7aFKsMFnuys4V6PXJrNu0tPkQFNwFoCHxFxROHqwZ
C2rS2E11Kc1dlf8gd8mr8ocq+C8zEhWQIV2M9OOCkx8t4dT01G4+sOEoX6rvBIoQj2W7pHGRjQuf
7O0eupEl0hFDLrsVCb5zN9oAzNfNmgr2CYYgl+xY5BKsRopObrxdK+a1elRjDqgEpyzCapERnBIP
Hi4Pxzn7QeIAMKchJ6FN/+LzyPG2M7SuPmnx2xZQ8UsIrdW6mqbe1mo1SsnYOPgkH7jIY+pyaL1q
Gb6XvIzbTjlxlHQNdXEwo91jSKiFWWcY2RUmq1rVeNxNcogJcxrpvMLSXbVeYMmotrUT9Llixbcz
BRDKPd9b1brcJ0dTgsIl/ITnOv6sxZbgEwtOlvIoKScUmlWq8snpyYRd20920IXU4BSKcjlMv7ok
xIZhCMqKR72zGoW5suhl5NeL5S/q7ZWRSZxPKjCZ7jziYi346iDKEHnrfgSD9Pi7yRUI59iIZmOz
67bGbNfpDlanMkI/ATbhYD0H8wUikdtzNzrOEEznT6fLi/KG1fuWCmIKlrYP5toD3xsi8oWge8hO
vgqMQVxTgCNujjgenr9WWeq8Cm7B3YimNWo3z7vYWQTS3dFi8ezucdJa6BETM3bfKge+KkoPHJzX
0hYsAS0/YRbC9DyiUqDkgWOgI8n22zC3YeZaeWHWnD4GNxRQyhtEuxRNM1nLsRP1mWOlZQn/D9kq
7Gc+b/AutCN5MpdfmNXXr0LdLJfByDDvgqdrfJVSzsw1xs7zkY7GKFXlHLl2fkS7dEeXxHpTPr52
+juj9rR3jWqccDl+i6aEapDd2mDDk7TpONRRpvSLU7UU0iWhqqWuxuk29lTnXvU99MmTa2E4Uck6
0YNRTT+Iv9GGCkQGiisUYnrH66PT0QNhsYk7Gq8JHKoP1e3DGo9Vf8ftAd9CiEs8imQ8c0Bk1HvM
Sn25/3oBwa+NjFRh5keihI3caKHDpVxWWYXR42vqit/qVkXD01aBomjsc1urY1fHXQm7ddwEIMIR
BQehDPzx3RSMJ4xJx/gFd4zPhAi4qxb/ZX5VrxjsvQ1b3MGLNnbyHsDTrfrPj9W/u4zHXYS+30f5
P3fGc/oSsb89IFA4+3LMF5jUdTHi7h8OWjvx8PI3QdNB3iCcdwFfjajZ+ae7KhpdaBNq6Q8Vbirg
1/CFBKYP9wlnZBpVbQvhbtAk3fEVvVgC5sbKhXyv38f2TcWDXVHV/JZMW9hkWYsumU+yZI3bWP0F
afRDh+xBoFZtKfF9YW7MVJRi/bI/+CiDHAQk1Qyp5BZumVDpyHH26vwfDFgPsmvwWlpMwjZzVSxB
AWhzJfJSgZ5SDh70akiA7WlsZJeXvAERZzBq22eBL+a8Zc1jn1zttTdpXJqgquZ6GLp0NJkNnP6r
gdfxcrZEWI7BI70yhGYZTbJMKZj1bB80/O0e/jfOroSiLHPCqeIS5f/d4szIzWRS1HFHRXFklyKp
qhebc8CJuDmZaOrTcKtlL4P25Quhy8MqgMi740f+QWNvnJSrtgSDhvqIHnd4kFJzaSdEdDeGCnLs
PsSxQhP4r2KjjIUYwC3pIkHStY0LzkvKtqu8WTvyxc9TLQRcrLuOYSPNb6/xV+QQWOEDX9vYpEQC
0HmFwUvilTqA/hg+zB4yJ+oeJSQG9LVsbMwxEUChA2ZNQakj22graMjj+YGhL7QtWkgnCZAVxukJ
iBvTbvxwFsD0E8VeNLrXGNy+evlE9ywEiSpqKe0Eg6VIFdI8o/+37wncJHNGqrX/Bh5JwwRc4m7x
pW7s1wrwkfZpeCBJOua9avye+uhCJPhBevgXzL04N2/u2y7B5kOSfg0mrw3+SJzpBaLRYwxXztU5
gUDiDUVsXn6PUjr9wTaUDYIGJV0JD5WR2VRMnJXnDn+w2fqvlNb2uAJJiXtz9p8AlAbIjN78yZHm
rqRDk/Vg73estziUxLgf7CXUqw7rNie9MleIEjvtPjE1/lR+J4SbjtrfGzHFdza91LTs1CQo26GB
r3YY0n5rq6UujwaBgqhJgeh11UEuItODKoUv0MRzT6TPOjZzvt72UvPSZD7kMLzAosvNdwBsxMys
KtHa4po9Jt//bnoOr/78tWiSbCoIdXKc6XmOkU91NNtzjHxq5i77xjYscq30WMkUCXOU+269Yyrg
I8Tg8QO66JVJlQgwku/oYPdPogvvVyDAJ7cQHCMklhAX5FTL5UQB37LTaEAbAs4S8QI+tFFeIkkK
F4Dj06OKXPveUQTVlMZakzLzp9fLjForyi1erY5shaAs+PBGwnRKXWhT7AW6/MZ8m3vOdjd61pA7
t73QtXx7HvuyMXJhfImkBX8qh5rB9fyfWnEfl8r1PS7P4Ztk4f20jqCoqsUtIDiXuoyYWPwWnDuc
icfS55ewl6Hj4XAG1TKzZd71YyaNzUfxmGYcTQUqe2OmMPl7rxfJXUjzOlojOCxM+rdeDcbIkXkK
RbFndrnpQlvqKS/Jo2ZChPMgcNijq8wvYeIe1x1n+hBQZe+CU2lRSxfcV6ReDRrtOxoRO1bIueCn
BWel88F6DqFuS9oZSOWPwPCa3jIt3FoikPHg5jL7LH7KZFwBX5F4RLZAFQnZq/Kg090RGSZe0AfV
wKvzguKEqIVbwkQLIOioNPYM1ZiYf2W3JmKIbF1ZjshrZjH61QMGYUJ+KE8JCisjfWK2tj0bFros
g3voSv5cEExCcxcsmhdOIfge0rxJBucbBLfhZdvPWi17McEEZ5WtF+dd7exxVMrrsngCge++EniS
CVnZFkfli3SA0Dvy6OjgRIfUud0S6OjRYUmki233mtd8zH3B7r47ILAtCHdtBQU8rHcEyvzQoFeY
D2jWToRRb5+/zceNd0MTWEgqNyMp6F21otxx6fDwaERaYAEy2UXqv2xGyGyPsq1FdffWJMlIzoNk
wVqD7CedP+GZIdv+aPLLjjb2C7q6kxP91r/RsHNPPHqWks5fGpSWtY9sQKD5emVKAaQ+9kKLF62s
lxjH8sCC3XukcYOPuN9Ez4iI6EDeWDkeN4rHvXSz+El74zuojMyQSE8a2ondhQAy4vh6fcuWTJEK
NBqsAIs+kQheyfcLobG//z1GgVMbP8aBM0AHlCjTk8XyjIBx77Rr7ilElQHrLS0ZDYg7MJgmOLSL
82Wmp1KJXYAIsPZiMCFsLirBiTk9OK49XhVX5PF5mtImYcSyY8meQ/Ms8w87eU8tNAaxXd7B/oq9
T8556lA3VXf1frA/IzdcZOGphYwbTne2mxaoXVAb7clNL61PWa9VtiBtLMiVBQKhUxgajmyKJ1ci
F2p5QnPO6QB7C+HppQhe+VxfpfsLYu1hUlbtI+Cdm+CUD3u+4qXKY73cdZZ+bFgOAa9CTJEHNCMZ
E9AQybZ/V8j55dtiaxHUUq/K/7eDCqyR3C74DeroH1xef6M9BUzI/LhznYzBSorHzOmA8LY5jlaa
rRX5BNlgGp/pPhWvxbQ81O5C7oo5sjrvkRDlF2md9dWFBBDGOpmIRI9pIArXulw08qSJ+s9h4wQA
RlrQwVpals1oJpIsprzzq4TAxGYgZN/wix67JupOEuVl37hr5vUbP37J5omlxAHeLAnjhaXwTv76
kVL/6f5vLRaNyng4CEOx+94xfF2ETjzVHWvljifn8etM6xVHf+BCQp1sPSwpcoNOJBeDibeP7i1j
OsXu3bspMOJH4rXOPjlxnt7zLJcZXHXQsmaZTPDtjzlkkEX5qzFb6Je5aJMP8T7nW3NIBnxVvC3j
Y+mz9kMvcK3Lq+CE7+yvcpOoo9pRhTZgLiLdjTZBV91zft7PZy41F/ShOH6KPySwL+mDn9+admg2
QdxhO88gaz7PxJgFKuZERBRdbk7r4UyTaKW5Nu+dKI1h0eBiGpVCgLxQ12JnHWqvSgE2LjLCXgQq
nNDZmxk+zwoEgVYWv0Ag2BFwYVatx8ic1hmKggItvsgfnc5QiRtUkCpty4zMYYPWZ4pg6GxryBpw
tq11P6KZweQ1oZcSvCJrdpOc/JJ1VwilKKS7ViLiK/IIAURcnlDB2qoasIL3eJdKqFrCS9aYWhKb
UMiw/THbx6WUC4iUPPLcDVUHxkwpv11BIHzjpDm7fh7uwe1KcKw6g2L6rf0nNp00cRH57VsDZ4zY
74POkTkRSlUQP86EzeE8wbYjrMfOEjEqAd/toXX5LziQ3X462Un+6j+4Eg0Hf83TLBG5CGZK2R6T
bQLrPYbZN6o2mGlfmKqPLJh102Q7P4up11IePXt6MbXqnD4QskzAl2QTQEWRyPyv9awkuYGbgflO
uryc9Z5bx/S98myaBsp5dFywWJzJdv85ehX/oACnD8TQw2/rvBCOW1n+QXmFKvZ2gtYaW4UM9yHy
qsM+toPFFxSGzWPyZssNyPRg4C1SiHtRopgcheaJ/ukeTQnDvuNqdesWnyRmjPqZ/ifShr+dTvu0
6erTzbtvnFvP9cU7KNzFB3asQUSO40CblrUt+ID8935ABsxLIAqTlJzCXmoqUVLCweNmibze7K2E
9d2HJNOd7u4OyhWEfuApa770GxK9gFaRvb0xyM72FPFrDNj0zVNW4jt9Cf31KCr6JGZfc3a92lbt
2S71vGpdoap5P7cLYj0nUQu6R1hgL97eqODBRbuQgm+grai3I4/iMtKJMhiEQQBq0GZKx18zCLQP
zrhy3VmTXHMKNsMzXxhCBbc6gMvv2zbROzmw6orH5O4kk+Pw4Yrb5bNyVjWUqW8qX/QE/kf2wzvN
ujEzZqIDRvkiUPUkI/lcJsQOGpW6cZoo491T2FJ05d+KFM7ZTQMhJJWlsrso626mG2n4QhJ2YL3h
YampmYZUSTpQsVezpj+55L1p1AXRJjMhAVZQ0YcJ3lUVwpT/FpOIM537bmz2ytzJcE32vDdiL8at
zMl7af3tdUz1AnUsr++3sWWXiOjrXIvsvU+pkmLT19PYJjSFHfSPk/JIi1A3sRevW1m448XR1jQC
8Oh6Zr5i8RPJUobO5GrEKK1PcAUDBg16a7LuyXuWXlFY6Qj9n4Apac7ilXoPINkl762oSoBFGfBO
cCW2yB+B/s0Cu76K2Qq8scPg473HVlhcD0j0nUg0Av2Mo6iiDnlsDUoe1eX8045E/LDEzFczC50w
72q5YPj9siAkybIdCcv1aPDKfHZnAp9ckkSEGeuXt0Q9v8PY6jRP9rqHVcVHz1R7Pt1lR7yHBryq
PVbNk9JngKeR36KIguO5bOBp1n85csMst5IeqAmSyPOtVAjqQsU+1okN80eZSBrGQxL1JYWPy7VD
HGRNoebEeSGVGatNWGuAs4u5v9ufGTVg9IdzvoFgJkgrEN7EINtYpxPa9wVu7DGn1zpofTjx7YJw
1jeZMgZokm8KPRnVLK/kNoaNTWxsB0wmCF1evA+OvUiImT81ZAQEc+Mzurms69F0SdymVRjKIv5+
H0g93P4P0ASELSY8EWJ79LmCiRkEfen/nzGehVJryc3roAj/ojy1c1OL1roO0nRweawuVhZ8PQxZ
OyhVHgFXjLGIBfDMLrMM0Y6+Gg7wKRL87aIWNcZd8HgXlM8WVRdUL02SiMVHvZ1lg7pmAsYOcSG3
RT87dZXCXYGBM4GxlJSXY7ja2Sro2R4t6Ch4+jNJXo6EacWSjjiwmzhsnGE8p5TC1ADTcpXcRDGH
5dIMjf1RT3TUDzAOo77wejX/qjLIB8lQBbkPpz5tvqvTQSGcRywK1f0IQk1+B4s8zQD/+kcNg8rV
NSASMqUhZNy0b7fodxMkXBYkpLKbfEhFuE/Z0KRE9RIElqAA0KEzjm6VFtTsdyEE7jQaWFKU/ANb
ThAQj0MpcguWe+f3wgcX5jwCmUhDlArUS9YSaW3qRQVZMwU83Fq39lQlAlXr23DeN6mAPrDoqnAr
ClW9JXsf7sqEgPEHm7oGxS0zcmfJ/9ZGLOfWnQQndB20BumsSsrRGp4mHEDzFwWLQH5molYS7id1
ZA0iGc89wifBNC4vCr6N3W2oSvlZlk0A3C8IBCd/7xkSuHSxEA4IiBbpW6Xkg1+4ngCN0vC97l5j
mM4VF7PERH2WJbaFgRqxCIJkqNWy5Eit/x41xWTEWiJAcE/R3yWi3yKItqTeY1/+/9UX1lKAuCEh
cqF5+PtpwgxO20Rqf6DanEQsW9KcUrYj0yTYDYQTXyjjbOy4uRRXbi4ED8uw6FaY8i4lfB3efp2G
zx8aIVbrhLeXmzxuQgSkNMZJqoziSJhbDX4K90NfhVYfTBGx3+BIIasJKHistjfztNXk72pxzbqp
TSW6AH72SyBtfq7dwin9bZ/d5xGOCX3J9FPhjddp4nIJu5+MH+eE15OMuEhXW+w4bjqZePsCd8mh
hxexY1E/mCWC61T/qpD3t81E3MMpJ0phlBq0apPqLUQTVnNyrwL/KXVDqtqAkBTGbWI9TsIxzABE
IHWoEaFjEdFIIqrNiiydX/DNgPJI+DuYQiR+D1LqG69HDHj72We9MiYnK6o+NNa4/yb3dmyNejDG
ExgjuC08zbo2YyoxQFsSPRX6nUROY7hFAl7CgiFFKOnZfG9P3G03DFZiC/Qvtdq578oKfh1K68Rg
SAF/4a3cTsie9msvDjR08XDt1dGaaZXPlLV15v4t2VfGshPgfBLikGC+9y6YLX2+KxyPRo3Gg+yd
4P6wbHseQZezN20+3YH87/75MuBFnXNE6Oig3lglcLy0D8/8KLdwu8kZ/Z5sC+eCL4jZR3qLj+KC
aWK6ZxvaW77WAlVRaFiZLVdSUNscUpXJ7D4tEAdeooc/Dln2p8DcVmflmsTImT6QnKzb+qliNS9P
gvEOEbCZP7erHWl1dh6IA6fMXFtOKD40MxcGadmG+HZRa6AvdKSL0vFDoeYn4NBeE8lCyXipF1Mj
FGWenJKjuZza/1sTb+QnYADl+5Q4m7KpsK8b4CW78Y1DX1JVUQAb1IP8o3e0pO7e6yz1gOEfHdZZ
eDWTSx5ue8S633l3Sh6HcxKOphYtYBqw1hBoiXBMOcFVPR72Qrd7eHzdGtrkb2VJXRWaGUvPQhj1
LbolvmcyuYk0c0kRG6FW3qFzzFO1U5pQ5QtsuM9ajNbyNnILFOLxqEt/6PMCKZyFMnb4iJoo4FfP
E1AEqfMyBBn1EXJ8PpWOWybRR9acMH088GE0kiULwTzS7VU/OUXSNCa+kzrROv9ba3nnHd9nBGu2
TvoP8wzY7DUk5mfEsxTIqo9q/Bg5bDYTg02BIicliPV/H/PM5IGAelT/bYnvNtVW5LudzgaVbe8H
pZb7ZP/I1r38AoJM0KmL/d4sW2KR5mzhEXvFjNtLuC5R2T3T8zyo0E+FHgyRb76Hr1BroSMWYdKR
sbzf4ynieq5mwsu5dZhKFkUXVdKLjCqUt3fR8dqUpl7tmsV1TZ1QQLJwtzIrUJEIWDJVR0X82e53
74Yx28vommEzg76fA/F4Yt1r/KV934d12oscExY/d9lqgqvpaPqbsZnOPj5dnn313XVXZZym6dwt
ZhqFfGE3/nbszzZIL9Od+In3Zha7UDC9df55W3cCJ0wkNrQ+tjWnIzWvKM/B308TX4IIENJCHDND
8vfK3Idtd0+gMf4W+VFGo7S2OgeNofwEkUNpW4YaO0phY18IpLdLL/wCXrwVU/CtFHNZ80IiCJsE
fgxydqCLA80XfRXYTKsBy+9wodcupkMjmh7DG2FI7c3Qa35LB7fWTb4VaaOl+ArKJH97w3WcdFUU
ZHouFdQuOAY0MYsjt4ijwSuDrv/LUE7SIU0HZtPqjltjL6FktNvcynjY4BdJu2nh7s+kxoBXhoQP
Onu7ZM3CzDdiC/dRMUPC0gEUW7dMD2CY700OezmbpXLjagwIJBuQf9m+J/QBwCFrghEe6j/wAWPC
i+T8AqWrLMV7krNegkkDegOjzzB09cUgolZ9+xz9J818dwQGKixcRd2eJ2F4F3uIaUz3TopWnBAF
KgRSua409+FwmCD8E00qhWr1tKlG3T96uZoiEtHqXb0NzZI7Eaw3vmdlAjkrmekhWLiMS6e55cXj
Xue3E0th1huj4iVI68+DpKQc8lbLyLqbVLW1yJVK+HyFNE5YIzgexeXohtCZmxwz5V6h2OVicyBc
BYZI9yan9H6tYEpjd8ryfGkpt01EYQ1Es1zzabJshDQHh8c/pMNzdgdZOq9xoaj3HiC0+BGP2gXm
P0mYKX1n184q29BJZ8ch+Qimjk7nBCl3mgUurx9Gc3s/EdzIznB7DacyzrrBDyZYnK/VE6Zb85Jk
lcLt9QAiaG3XXpQnQFXA3JTOzasd+M9hH/0xcwTlENu2apcIJNobisUN+ki2jacO+/a/yby9GiJA
hPAeXz6lkFAWMmmfaB5+0KW9W3iL6Sx7jstfnN7k8UO3ngL/h1aFK9gzPfCwuvN6P9r89ZsTfV4X
l+EOjIo147NnPgmpln4izeknSdS9rQN60qw+NAVoHyG3gmGe5QMrzadbYJPI6bzJl/r7z6Q+k4t5
O1owA0qpAAV8OmQ5ncFqFHzRg5kAZvDfhWVDNS+wa9f6Bfad1HkFyHe/PFpvCwGJr5QkJvYF95O5
Yd5qTJSAtnW06kb46CCUL2qFNPEXw603vnE6j+RgRABFktIzdYwQIGjk9lrjFGKpP/DwwBKKkqbR
37abPkKgt+FdljQXrAiWE0Zt+JXHPCHlOKUo/uPIdTnJB2JDDnY/Hp8S5R/zo0cDj0WCLd4tWCjG
++7/EfZ0hsJmY7/F62AOnrzmuIys0OHFxHjSDGlystKAVimvoJ2L/hf3ygMrVLep8fi/z1TUrOn5
JyBiyCt2xrVQcVeUJpsQMrXCzzarg8n4936Ctd4Bw6os13O0nsQft5bjaGPorRlOigReAPWOSN/l
8uz5CANjkxJLvqavvVPVzfCd3VtW7OXFU9k2fYEfzzBGBg6tS4s8ShQfjMj+sA50Zk5v2eGogEFy
wmF293fdCYKm9RzPrv3M8PjEoTmHxkBONPyVg8ctZb/1iPmAWnbkPpFKkZS+Z/M44rTDYVvn7Vcy
Tmz1N7s1I87dpEJoWanwzAOK/YVBgiIPvup+d+oWJE8Jsw0Dhi7L5kpWyLRJVWdL9nh4Axtxd4mT
ewQwKOqeMvfWCdJlHlVeYSuq9Ywd9CjKuYKONQgfO4vlodL63XTuv+QihfLI9+ODU1gZ1+cshSee
FEXFVWUxJeWCq/X66L7FwENCVFJreUVfAq3uik88dBpHKzC1u0PnUGTkfN3i1cTUmvWIo8yo5e9n
iju3Bc0HVtCVlBletfSFr6EUc69DICyFxC0bgHKMRfdahdl17C2qyfiTIjkzlt4Qx0ZBexr72mOo
Ta83hqK3qyryxbgLqriQhF8j2cxpusYxgqYewPob5YkJWQhw3bxRnH35P8Tm9lvw2q2/3IqSwhW1
d3Bp0jPDQm80mX8UhVvna0WUsIjaO4NTD8O7TcxBrDn5NYwYodhfXetDsc8ViXvKoaZo9TuD+7Uj
gMlHjMarYPj+iNIqtZ5A/JzF3A3GW/kHwDkGH/LKsbI8ZkqhYExiyfeI4zvncYQP++cly3j+oVYQ
wDDhKFwK+9XKuBxyQK9d57TpIS0u1Lu+N2FNHIPRmgu75jpziWBuqDbL1q11V7XwGu22SYMrgS2A
xVN5UQp/LmAVqVneGW8zBdJUx8nz09UbmJmPN/+iivC1dTIHs1BgDlVw7qzOAPAw7FFonzin0SkX
ZzbQgSxGhWQanmFxT1RApZbNzGjiX1p4zFi94Zip9D0IIHfNtIsIfPscwmku4Yoyy486W2LFc1Qe
lrqZLPPo2xR+IhusgPDH0f+azpoDmcm5evl9cAX5jethpgqjkOBE6zZKpGwa8VCO929rmxASoVkI
9zwSlDaeh5jDBs5dG6UCtHc41EFccJL+qbTX5tN4dbLYVP7N4dKenvGO8OBCgaBtP5BW0PCz7E6U
wLLgCrGaXrkIkAqpZI5VBZi0Q2tz1XAt27foiZ2qZuuyi6SoexPLuibvf6RCsUTVBOLL46tVvMZE
cW+pj0wkw4VQnKIE914zd+k262Q22A+7jZbDBFUiPIozLL44yfUZqiX5aZyGGmMOpL+a6R/QCkZz
0Tu5j6lVD7Zjc4BoWf0mUvF9WquoHQkeddwiU7bud6/B22ZwwYNDJ/DPP21hQZccrv4sWzRBLFV/
ktFVCBrpeicG3CDfkZA2KpSndb8TouqNZG365OGuWNHBIKjiyBGG+v4EaXOMPpyRzAz0JcpeQ/B0
jzf8jh7w4E/RBtUYxeUrBQvRZnHIpWmlpZYXgPouW3rWMvOIiBWpMzn1gGUpkIIGLMaWoyE3jmS1
MRLqBX6pGXaH9fVD0hXAjxeX9M/RK5EDL1ANfhq1WGnYZRKPgwvyW8YMdO111MBVv+EhnE16u9DG
L5PEwQLW4a6ysIbw0vsGY6kLTaDkDkRN9nZRZdN37qVnOoA9JsiKVv/1l/4+qNQVYVaoJ7G1dQ6K
BfTxK6EzdOyU/AUGr1GBsM6vrEpVRzUbVjo9lCKdA1QgWHTSArpWUWfXbu4uDnP4wNGLa6J3dUi8
nhWaAIu9F2T0JdPlQIsCHTeSTRCrWzBMovOYUbNC/IoEaAuTDbsKiixbSHLdRQNkQu5dIr8z+jbq
+xnBEtCCTcjd4QhsPRIHiZC70MwJ0stmWKgXsWhJWQRQJghH6OnB2AQe5KXGIPeWSZp1RVz3Klph
gJBM137yv8qmz1Tio7WeFHZZTLw0ObuJYpBqWGw1p2d/6fWBkdrnQedpUWvUoWooc+95Gz7K923y
Du0kpPRB7d8GEJfhYu+MufWWtR12KA783MSJuk3v6X86tIjG1ce8Ta1jJ8KiqttHACxDyNW2mUil
9etHul1bILs/tkqI1UuQyyGMQanPtxMK/BFBE9nACZvNtE+XMDII21xPcS2BpwFjNl4pJ5FfcwNo
nEunG3Zwspk1tLzR+x7sAZOTkta/2IJSCOePH+GBbznjlYL2oXkUeKG4OXVYyGjxsjfN97ZqwbNm
AJYgbkSp1dPC4B40or5A5dAu81L9+FMk9ctyFbTdOzRuq6DGJGWHoh1e/dBfhG1XatuZ2eKREdJ2
GQ6Dr3ywRj9ZCujq3uaoVwQvisuaDeLXRKJ8EV4sgMW4+LTji6bL5hMVAILSHfgDykcRiuTwugcJ
4fe5fz8i9MBqVIuONE1duxbPvYxWpb4dIhVBFk6VdxmW+HzmFgZTcwrQRZWuOclxgfcVy7LPyySN
WOL2fnEQrgIONS7COMubKMNp8NuHcFF9YEtFKcDGPHx7+IV+NownI/N59Y6OaGM9FKvTwGJfWSBG
HWUdx9qp83IfRMN6dm7DHDhDkhwsM4bjxCW6lMpgbWAAZQzZ+LUqzGDJBZi3nYLQitsiK8zm4Pj3
WaEyfxa4czIFDVAM4Ark4AvVIPXTL5L9egiXxKqEh3J6NbgSbSOmrFv2y0kSL23uU55wD0EnPjhW
2IB4Q+eJtBwQ8WIk5z/t9K+3ChRACpoO81QMIEeIqStPJm5BmuRLiGYbotoOq+EUAHHTWwT18zPp
1oRhLaZzrnHTy4t8rZ3k/WbBAOalbAgeu8pq2Dx3x2G0vjszU/Wb23dOzgtK8TueXzbHyrjNhui9
pYYEJMG552HaNIwB7Ny1nyCMEj/0DcUSbTXSXHsE5JDHaDL7JaYaFsB2DpEzZcaR6Sb8wxuUnknE
lSoIcyn93+IPuPZ5g2Gn7yNmaT5WBcCY11sGOzAOK5jhjRvOgpC+4kxXcbS/UZNBxuE8+EA2i6X9
MHOnfyZAFE4I4DwUQjq4MOagZ8xvTUjeA0bzCG+yXIfJqnxkmuXQxM08DiBud7lxAwX/hu7EZhda
MZxSwCArvex6B1YgWXDzdY8dXcEyTXyyiq47soUrdWaHYhFqJ7igkyQebfEODZ0A6hZcCpbdz6mj
GjOIpiKz++hMBCzwFZStXTpD1XmN2gC4TmxWvGCHoFRUlO0uuvyfVm2mTCpb4Vrb99AGeHcooGgz
EOgTc1FuBPAOyOzSFotrKiiIss96F4vAjf5g5V/GAgAcR2HrM/JKHByLRtBoZbEteGBB9B4aDHin
4/iwKuscW88el+ihucEv0TjlIR3cWCrc471eVzQYgWQWUMLNOO0CBlroAvnvLgdpsMC80X9XAy5J
g1vzHuAq0XdgggkEekgC0N8BSQDMGJIv2SxAK6iiOIriTjPefS9RKbR24TnRtI0oFIV/ZEuB5CFS
UUUM1Q10gfl40rdRFnb32PEtF5ho1sZyRsS9bhEPWTI4dTyWpmJwQNUlVaGw4nZeECLuPluEm0Hz
/ngMlQRmp4/OddL8ddMUL/nr0cjEewa8+NSrxQ8PQYbZenqyWMDGHN1F6GwQFwK9twki4KUEOwHY
+RE5QuCI4HUyn3MzAcY0Pqufy2OYVkPYzub9lXUAaOj59YibTuQvqhehlkfbju7l0WVJvay76+aL
eeHdV+8I5/bNWgHfAmREFusOsaa1YnkHMV7IoB2trpJAV+Plnq7J1wt5AvQBtRUnoIRX9tjGMwVa
GsNFAEkGvtiy39wCgSnMf2Dpy3/DYtncwZikiyqFWAKNe3xx6LTP2MaT22gV4RGuBrxv/aSFRzXz
kiuMh26CZ9yuGRc9OV4yh73a/q5MX1KqI1NgdKzjfgEANbupsNbaCdZDiNQyyJrYzQED6bg5fAOu
/Zzc59uaVBiA/7Cj+pZmMa9TriZMny724sMtbB1OPKudrxPOCngLit6pgWyn61KzfC8pncxZjNI3
YcGLgeVsxKpJG4sY1iXAiPF/x3PVvPCbOCjQw5n5AWIKgOKOjDIw8k6MJZQq5naFpHmX3M0nlsvp
mcv2ehmzNXuBNiAlq4lh4KbfRzEoLlx1WrxWEtF/0jWq8zbflurZMRyXGmHK7CnjK5aVV/rAnY+b
obliwidiBCEsnv8Y9d8VBvJAc60zc7HevwMh+aLPJsSf/ysIuoS5ewECGQCj+LP2/kgpo1xYX2eK
vRFQNZrsIjhtQYNdqk+2WuywBgZwuPn59rfLS+ztv0DL/YH4gbTJNJRQrXcogEh8sOyodCN07eEP
57oplMfbk3cPDdg4tJj336P9758GZpkEKQl8zzq4JGiTn2n4gwmsYyd4zq+HsFH24L4OOap5mq6Z
ZqwQivk5jfAFbOhUWYsfGH2BNN0JA/omNp1y2nIKF69Au5oNAse4eGy6DXji0SH4isdcft4sPQK8
7iM/utpbkRnBcIAx6cqA+LH1GrCYKeHqa8Xf1NK8Ro4z404QvT3ev5CHz54exmZbFmXef+G+vuMO
nw7uBxBcIyeFyrebhHbz49rnhi6ShL4qz4i/rTUear/ANRL/BnE58VL9jhP7kdwM95cXwUQm7frc
ju0EHJ6JAxB6JrvKo46E72LD9E7Nl6nkbw0+Sf3644Qw6JKpVYZlHx7SJhQAiYO1gLeMbbF+7sRQ
7qnqexE4ysSNjvKhBcu7ZRS5RMYhlmV2klVwgK5I/AgcgagaahJKJzQUEHfm2DN7e3mVp+71LwLO
dPZwAqeZDGQ3AY7q/xfTawXXkavyWQsVJ/tLZ8cDOr1yDbSnlxPzU6/RQ3R1EngyiPvEGojmp5nu
z/He+kQTDjsABYmXzFJ1XwHM5pE7tVxez1VCFsXt6y1FtK3jMEAXY87L1GlVWzc6sbC1r+KowkDq
SkNwhFGkhHVak95raJc49BUhKZjwBviWitsX/a4uu6JAi74Lja38UPOhzUvMF08/mEX6KzdYie/q
L9s5C66wK2UNwKDjRdrEwvM7Fm/WBGha0tDyXTfUbo6tzd3jpngUOspOt+oKijeqpRbMJ0HZMZyp
05MsxJ4QKI/+dZ3X7RhhzdXUUzVHhNWoWbPG5RkZzfCno5LpZykPMD2iLBRT6OLKcWchSVvq4kUo
gPkNYCvWkMjyG2UsPyfi9l54cwm+8ep21hCEU18am+LmFyl3TcO19ftDAJOJjC7jpLqiwL57zpAd
5vu/WqTntcKpi6p1bD7NS7gEHw2LCVCxMPBosya/XKPLOyeQ1MYNSPy5C+MinGZ9/dWDqjxhebny
5U8DwtuN8k1Wr2VF5LPnF2e41/ghrmh1CP+U+RIT1ZKX5H9J/QpBHHRYUvjmR4ZlzU5Ip6Pj1PaM
owXB0oEwwhBfPKJTLo81OJ0Q0K2mNNpJIL8F3lNWjv+S15UAG/GM32DHXsBoq+B1n8SxEsu/KFe/
2164M068mylEWGLyZEl2wppKuvzsiaSbCcXn+ZV14ucXFK5HLRkzZNnIeDh19YiY5/f7yFPPcyjh
XbHJu4AL8VixRKiD3VIydIaTbn4Je5cP1xJxtdyWpkipc5lsLrYOm0N7HtZKCF6Vjhj5rr9oDb5S
/gmzEbA+1ZIz1lM/+MR2n1I9LzTaF0Bd1kEL3qIBfXekLHHmSGIMCeCx3PWDQUiqtOn3S0CJOBn8
p9S+BBS+jRjU9d/kPSACXUy13KYzNnz9n9myqDB0ShspEull9ERJbJF5WOgYJuIvFKguNn//NyLa
NEzIB+dnxuMihsmvIfUK9ENUq7k+oxalfRa8o9Nt2zUyZVp2lVKG9uKwoNin6bayTR13amkiTA8W
WYscOF2OTQtUMgLJ/+au0zPn1KRvxEVMoSPhKqEbYW/291Fsiil0DzL/LmhipG6fySpYTNoxvavr
0xa/SeS3RIsxvqyem+lLo0hGCLj83gmmR0070J8BPOc3jVOO2iUahTmORuiNsTGRMz4Mir4OBRuW
oT8cz+nVL0RBOTrF4sNvXkoern/rFkbwkrG0kSHOb0RzBd1kNjCbuPDSid9h17gBd95FmkdobvLs
MnFfCmJzh42wqtcjIUlTV9T2rMvvcQoS6PFdyHf8uDvQIhcKGt+NkT6uPz3IcPSxPb8ycuaOzY+W
DOlkzuJUi17fSTlZJSPdjzLYpi11rLStFOIUBSVFipWwn+HZLXRGtd4PuEJphttpfRKq4UCpLlv9
bJXCnr3BzdFIFzWUIW2VT4/xrfiB9jiZhGRD00o0efvhIt2gJRP38FRJfrYz2CdUa1WEmJR5fzs8
+OfBkGvoVRgGnejueDlkdGnFs9k1orYS1GycAKpCoRUqqX3a7oLWVuv/iMBSuD8xDqqMXZBXv4sl
/uBVQnYCKLg57WJqnZTfASk3Y7naMIqtgGmh4Vy13RKoj0cgH22ts35HfmmVzkSw8Xr4N9miFgWc
P5E19MuFgaF7DnXapRScnBUhedxO0WS/2+Jcs5XuykH1tiTLZyTWKcs+DTWNQeCntMmZTWTxYEyu
HW4uqAaNMTkXjGnWdHgiHlh40AooY4lzSaO2TUVmaXY8H3I8HPSl0UfqBznoDkixJOUTJ3PhyFjR
ZM4KQ8+Y0RoXjr2FjhJ6gqL+GeKs+9tuRhE+Hsz2/nK1/MWRdRYt/nD4xnGUE/n74L6VqIKlZcaf
VhkKiMSKlDiBCrKnTSZaq/ppGew4ixcs4+avdwaeEvpBq9pmwKNn7GG0zmbJdzq2nGORWZB919cH
AvB8kkDx+KWC5fkUBQ4yoCwLHo1T2TSlN8KMQ2HQsagKCzEz9F97ybYBLTf1TXzi3dEzPdic/M9N
8xllhDLouEJVKYinXz1uiNeXD8JYXP5PBhMHJ2K/F7m2yJRsMe0MbvUMlQEqxOPeSAaRWKLLRBZp
nR+6aoGqn/CWXtRXPM+y2hXmFYK2p6TYpB1csCS9bAx3VL9CUy17zLPQkIjkKE4n9RobdiLvyRHg
AJVFuUXQvIrzdDh3or0X4xlZZaSZpvEQ7aWa2Z79u754Fjj9gsjQj7sitPz34qOMTmcWR+5wSjdi
o/UcakY7WiLyPHlN4rh8hr1w5ZIyXarfuZ14rlGsRZxg3yBkGRI8r3buOoKHB2fD7eo+L4NYK1N5
PLuBzQ//RXlp4y7GgyFq1io/6cpmt4DCPtHXXgz5FyX2miIUchqWjhMZsGfhVogr9KPef28mJy/G
l+NWa3T32PbWYNtE6nKSWd4RwrYF8RI3qwfAicAe4YYVJmO+v88db8D5mKwvMLuS2NsD1bDpj6DZ
XuK29yJc7/bKW3iITb4CKFiIQXthoUUkDDPmZ1+Psw5cUOwaGmBa9JaWU+jiMgHMzngB2jyvIxAl
n+yO/D0L0EciEY190bfl6CBwylltiQXFPRIDJL/S2AmA2uLoLiTzlzKHDgXPHy/9iPvsnOvvAWdh
CnOjdFDDp1x5Rs6qBXoZdFkQFhGDMK5WUpI/9urT5f4ELNRStJ/gTqlbeS/p1/zKdnUkOgbI4GH7
GP7Ul7x3BA7xrUgdHOXGhsbIPonriF22EH5jvlwoQagGiFyTq7HA3e9XdR01CXc9vnUTx+h3oo9m
5muHZ2fTqC8p2BHddLor1hKyNWZJDdZjjgHH1LT0xfLzAdzDak7GR+3L37da8em2FG6EXOmjniCy
CirPeRc0V1qlK+AFCd5dgIFBfscbNWMwuEFaAyQIIHuY3aS5dilbpA9+2WnsrSPYpbwi0qSCF32Y
44maZDhzW2CyfiiQXwzOLskVm/ydtX+ZjnChPE6ZqRdtmfSsdn1IJ2bY4GyK8i+sE6wmMcw6hO6G
ICErFtAkKJ6DrC75UVhUqTJgJtspRccMWQe+6xmNSG+ggMr2y5KRaG+MLMo54L15PIdtzq7pAPpO
FTtQbIJAz6hPuTqUmi9QsoFs63AH8wzjJ8S04l5DSNAGKs9okWi/niVkt3VeZ/oAQ12tkndsSeeM
/gf716JaQgOOpgtezKv+C0MYYtVmWhUel+V6v7WBBekOdMhct2zPwW+0CR+qTGHJHRl1zEgdcUZQ
LRYJD7BSOVLYYKFgnQXm/kdO204+gQKr9Q28AUUy4Xky4zKxsc2lYQSut4wBUrp4H4YqNNG8PJdg
kDeoccG55+1DQiiJCHMqS4jKnyQg9puBBJgiurv/YcyolMHhwwjNGUIPR+yVxgV5c6qlp+1cEKPP
317GKhtwAaqpqfNLVcaouX0WgG3jeOnhmHCPXkcx3WQ6HsRZDQeW+MaureweFkrKFCKc6O7n/Y78
rHA6Cs/pdKlW91BuSm9k84LUCyvKb2VpQJ7kXc84XacxQZBbeaYMCcspwFqDYLeJQBTBLarYrWJQ
TZcIJubBot1v5DmE1BBCGqhlIPseLKjUpefPBNbGncbJprNil4ldNuJBfp2GDI8a/lCDybDNu8w4
rw3/kRN/JVlw6GXy6tkgF7M8CRjb1u8X7IT5M7hnWR0CanXFBC+fifoE16J0T5/cHiVbDBgk9zkx
vHl3jCVQ2M3GeyJmkSazwMu0zCDoo5g/RgbbBq+kCbaq0sTFr5OvWi3kRo3BYJlLm/WyDdhLbi4/
gxMetfQ5i5kaVFCDypdz4I9pMXtOCLSb0MeWtoWG/DoA8PFO5UwBNBOFEbxVUTHRTeLgJ/CWghLF
iLJZd5CfWQ0zbmsUUMbXH6PthAubM1KST+aZ8gs0JSCEp74wnTZA7oT6TCpO7NzbEh9djHOcncZP
6e82VFBoZ4c8SuHEgCAqiBEHvV8YwjlVDBlEtFae6BNB8ICTaX1ZExkQpm4+Wq40hRogKlGq3c/V
BGOtsVjCvncXpPefdMP8RAKPefQFr5lZDOvwkuqpX9B3gq2y9lLgJ0N/AItYXobOHb2vcEnwF7zQ
Cy7BmXqlUc1tFFWGRJ6a0nHCa9FbqQdcE6kYYUEnXCKsw5q/BYEs00atx2n06dzdWK7bPsKsXq2V
d3g+aRBP2citsQ7OwyS6l4FVzfgvPQlq40CJgz8UfalTNS4Dpnb9GGUcMB6OBZnNcGGyvCqhzjt1
OAz/upVZzkIhn4F9k7rigjTqUqHovCbZA9+czIbxXJkwFQq9TRJXsdNrGGdw8xzc1D7uDGjMCN1X
AyfJTypRAePUDS0hGur1mRNBTTcVr55mU2XUdi/7oXfqmFWjQkRoGMsjN+7M7AHUwwcS0+JvOt1D
T1jvOHt8kHjXS+IKSXStQnA+1bVq+Hsa5qnjBEIUYq9JOzFn77DHQ0bfEAR4VgiUCOvYZsWgmTSO
vuisit/efOMo3lz1qxh1aeaI59EU9bXfk3zmu4g77GgH0Jyzor/DFC30mDiDhIPMSteloNfzNSy1
eYeEKsGOeEVm3NPAR4QJtImaf1QGlIOi6BLWrxClUSwBcKyTK0hubPO20pePCQOLNsVJ35oJHeU6
jW0dHHoDq/zCPGPPsnvSOMe2jooTUyJ9yBlFrHYV5rhcBBrbs7wc+P7ouJN2ndN4FXO5wcNLM/Fg
x6AYI1rrDEFCqtQyBUV0vmFXajKZ/OsZvZK2OScab21HXKjbCBZvjkVc3ZydZ8f9RbcB9x3dJiHF
UULY6M35KvVwTj8SD0hyDAhIRq8ifTwpuFyDJioBG1JnWhEgbpgheVeX0rL3I43yr6tki8bpO4ib
19v6DQC25fMAF1Hc0G5HRTMFU0iIOx4PnI98bcHiqwlXuSNJMoSN19q59OBONXqeqDEdRO+xTYHm
Lo3nV0Vtz0Q4u1HZWEe2yPqcvJNMHJYZn9J3ed5JLRlKPfbCSOwR39Vg08NO9FJhRcnpLiFwf0CL
I1/pcYed5EWiLuo94qPAQgUhLGTRndOG4mLgbekxW6CDIZsUT/PDnZYPBi8SYLDfyBk1/D+miqCM
tAiQmZXDPbkoHXsyNXPvbgfWM+EgKFgHxJ4MwdmO4runvGy2IT3kxkAv4v4VcoHZmN69rDiB0eUg
VC5ur8s8dxUCSANrYXdoj1Q1RH+Ynd8WuI4xiZ8mxcwLgp6DNqZWvcpGLHfl+eNPlYRjV9+GubJL
pDID3wvdBXCJ1ZaUT1q9USGy4EcItZepPAd7FkFUOSsCeIGut3i8j8Y/QgSorMgZ8oJ7aV9q7Igp
KpKtJanUOMQrvviofOY2GeSmeGsbZi6g7Vx0E3+mMxVpvRxFqYz4jDzhTAJATqvlebXJXl/hqkdZ
fYRdRuTXgyPrQuZKMrR46DU2Z5fy7rW3yNVHf8LofRyrp/bx74Bc+O2c1e+ljTff+27L28IGK7e4
+TrIgdNRf0tI7UeE9zhSHaKpiWd/ubKifuA032UjIAYgyXysOCmkIeNSFX4cFLgrm/maCsNdEBTQ
aFg0Nbn4ol94FALj8vDBUEy7iAG+j5J4v8tJ3zyWLTo0v6Jv4FHGoiWap5ryTkUGW2VZ5O0txquo
XYAdt2rHvt4G37WJ93eIIyj9T3Iyjz6xtdAb86/mJJ79KBSE2BN0CUOLVbkUHhav+f/XQwmD0oLI
onj3ehr11xo0o36AYArb1wH6gbY98I4VevrvV8oA66MMR/shCQ0ueR8uGuc5U99iHQ/mnoMFkU9S
m5oY+c7By1IP2W0GnGe3ZGrMOOP1qAWr0wjfIBXevzqEm4bLw1m9ByKVVRMVOPpuSFDcvgTZeRmO
C/2lloX/W6hqKwaj2XIezYTZQHIc9WTYBNam4N3bt3UemWtQE0GmOXYmY+Rw3zWosVx/fNN0mmn2
r22O4pvtVdwVYwKnRCYe7PoEm2kNuBr45+i0A08r7Rku1imm6xzbXdphBDMdKKd6NaOwdeo3Zk2S
5gSKahG7yAcKbfasnBpt9Y0VpuSeiS7TGBkF3x2KCIyJkwPiJtaVS3zjvnnjxbwsUVYJWjqVEA7y
6ipacRGvnwcVgoJcddgirTRdpAzRGE5tFYSNAThaCKwktzinm4//NvIJAcdO+tIqI2uo1S7F/BAm
9rQunmSmBhilWya0W0oeM9JJ6Hv07zzIOaXs8wk9J4nyUlxlciyLmZbTVwCzWJmmDsyCgZCaoFlw
GwZmB21c6ajbc+B6vummAs6nYcvGihZ/K6iLLOBPZcBhCwZCsUc8d3xKUVeiNfkHwEzNsgDAgIaQ
cr1ePRZrXSdjQE3N5/fJXaYjv3tUmpGbjDa2Ld9igKE1G2Vu1YC3AgZItuFG0YcDVKQaT5CZjVO2
YQDzSHDv37uO3UrlI0gSKdQPTxai0ATaX03XRt5sOz2hB+vA/mhInKeMYZqSVsnxw7Dm5lGUk+u+
ux6R8cllHR44PcUdHPIK3kTCkOZEW/auFnV44uPIYgg23iuKaohej7r7tMAPDkHEZJ3Bv6NNtND+
vTW3wwKKfLdhQjQzjcm4Tm4i5x1Y2wyCb7VwDJmPUN9S1LgabjXP9hMDrUtMBPPAFk9b89Bo4ieh
EACMBOd3MqTgldCvYVOL8BKp9dYZW+sLt7ibRzMk0LbdxqyrwKKs8x5QHZIpAsAGsggMfzkH3IEy
CxTJyalpwiqx5+ociHJj5fjb8Mkil7GYyAEh3yu/ADPUmmbHtthq5NEy+LQ0pdlj9gGndzorpJfn
iBmGGgDPi78Lbe3va2vkmw3K6d6Dtap4Avqt7dhADwBkjYf6pyIbLggAjCmSQGWxcCKp4QVhnAe/
c0rG3s2AsEMqRYsmI+OVPpd0WCiUdmpW1bGq0K4nwYr975bhxgAqYPjQRAbDCgWEcVaH/t9ocXKC
iRZo6ylIXncDTU4q3VRJH97wAoS5lKl/ldtJWcZBOUa+CdXO8EOvX+M3f3pAbau6pQ78vaCBNCL7
ETGFw32hjr3KNhVRWEIoB1FUtusxgo0LgRZXJpB62EVrJ/BkrbmCCVMuPfcoknGo7Mg27yyb9+YC
NLRXORwxx1W57PtwuF/F818eWOFXZ/FyzoSqpgusGsTDaGsUltQpqXB+UbDS4bJQsstjwLICad30
ANVkRwV0AVO9hMO4ep9TzA07BnjY+WJhRqIQXgClR0b2Gyse9sGPF4UUxAUFXsrNWEPzLYtRRpOK
26qa7nei2yzyzkZfDieYtVJfseR3k2TNcPgvccMKnyjjV7gJpVl9pF+ABiWHETum6bZa8gXhDse6
clvz84VfxeqTUXOcLIoGe2LSy1XJNS1lHQ8VNwC2tg0uYFKLl8CUCDqg4METa/UDVMsaWbUx/xLa
D8Asj98/wpFHZS75uHyWP+2ipWfVUrpBRMKaa5aPPyKizXbKWte4+wNGa6zSTrY+t+bnGp+gg+KV
3vN//G1v1g8wSmrCCExQ1Fdq9S/OWzvOlugyS91uHoByPbUImqEMVJjggKg8e+F0NTc2j3qftXYH
F3KGSfFwbJqRlIuCS6XRLL9v/y0EnRgW7U/3PpX7GAme9EDXQNqshaukyE/M4do4HEJzEzr0mfLX
HoAUp4rt1T12sp65kDm23gg7jPqc9+nI1yOGTSk9Rdr8tIClJnxyeQ1ympYEICWXTaBbkYifSN7m
5Uj9XF5Se0EWat5uazKLy4eKEx9Znd6D6yazSD1dqVZnglNh2hH8r5eOSxiOXeN7J0AIQL917rmG
DsZ7rmGJd1BmZmrZvebYDjaGlz39s9Z2qelyA7gEpyz/VmjCSXFw/G4nY2MQS9tY2xZ8Z5zwuO3/
cfKn7Xaz4vKTnqGyO+5790bA688i9wgpH0gY+NArSrQdtPA75yEe+Z06CbLoS30lNzItwlY8VDPv
lzabfjdHAC+HUPZ0ofoGK6fB+sIg6tRH2RT3yXFgB3g2YZ6+ftuIzkf0d9eLB6995GbahGQtL53W
SVAQEIX0JKsajLXuYeqHCbs5o05SSdbWhaqqaMmr+prxw3BoTt5NYILkHUoFK0BhY/Sgm5uFWK4j
aHkCHlyC7vijpUf4Q8zUDd6f4F/7fFpxjfrUvOXqY+wzIvNNZ8C4ybhGa9nYjgho25NjmebEaIbE
p/qCfayChx7OudkTpaojixWUZ4DCyaADuH+0g54CN6dTnCb6C101aTxCkKfLrQChSYiGnDPnzrbN
Ctcv+yW5keO9MghfRSUU2AYRLIxL5+Os01w2EejElkBP0kGmZjvYZTBvgjcz5mCXeeiQkqGTNa2C
6G4c9pamxXuDoZDdr9h3JJ6Kb9ZKoghK24Px/trv7yKpAk2nxTgYQUjRb4Hm06mwWFDY7u+G0iod
aGLzChiG7z6dBZU0wy9iifuITARpYxrDhTnJNxcs6m2bqNhfzsnOtTqs47uyAhwo2oKAWnwWx+LM
b9cmMeDGfFntXl1GmmLhwKy7t2NJ8J3Rc3UUrv4dTwt7hkXPgZeaLBxeBKWwHgUdPeaqK5ZZys9L
exnS0Q7c0zW0EDEm9TBYWyF/mzZvECGtNNgOHNPRh09EyioE45CFThQQqz4/mPnctvgg4h+Y09Fq
IiYpxvWjn41xwUfDkd6IBpltI6Id6AewQO2ElOJDh2CuhBbatgLU/YHvSGcevSFPe3/8gtHUf9iv
4x+GAdgeGE3KES6ya5S0z5R7a4cH+EPObtBx2p25zfgh+SGzkl5pDKq0a+uweB5zTuvKdVyx8VqU
O9UMyi6j/JGdWJbu3JN7+3qbJG8znMA1uOi4bsquckUlzFPeWfvkJtwATYe7wxVMXUXNT7koge5h
YSI3fOlAECbaiLeJMQ6Mr+iRCM+BE/9o46zZAA8srvAbUZ0ZeXaf7eOTyhUHXWMKVR4QrWwobrPI
dCtI7c+Oder7VaZP3OPEhDV0X3OAUeTYL1fBjk6bwgE4dKXrsz/2lqcvPxbAKke4T1fDp0Px73Tn
1lobOPWulGftoXFLa8ScNimbGfrbB/17gYYkWkfuOdZHR+EUODKF6XarJx6vkBRObJwuNOq67FIp
iS9r72HNbOdMqJbWCzqJth7tApFvsZiZ929ViNh+ajf2qk7dr4w/PPc2hAG4fKmXNv8DPsvDc3TX
1hjWMl6/vWz+F+x5mOsdU4N1KheWQ1OCf28DGIqJBqVm3CRe2O0SJgeyUNe/rUs0N3BiDrOEgF1U
Gv149LnkE1jUZAOxwXO9VhjB1ccVzNKLcny9FQpJeZLcj61bmH1k9ipWqgcRhahzijX3K7IxGvT5
yUFIJSK8QJeKQ5IHJx0jI+cESUE+oUT1PHWlziMpG+8exBpW8rJeXjF15hEYKyd3OJ870oA9V3w7
BwwI3jd4T4X23RQymxN4uKLh4b4/Zx5ALS6U3HEJ99+0/yAOzIYcGbdVFkhWf8sq3Wh8YVO1sEDh
zEBYH2YTRWJjHwUr4g0KaLsezUxQmHW5aOLOpfjAV2KyWawgnmB0dEQurHcnqG9HBQxPs+gafTlB
RFxgcRFkRyyVkaIO6SiTqVo5MQKgWHn9jiSNFYvbg1WIgxuHiUDLNMA8oS1Qa8agigKKsDEL/C7T
4hWTn81KAjCoAcdCeRAtSh74FoW8vpndVjrhe3NbJryY7H3KjKSxgZB6p5Ycn0qpSdr2L1sjsR5r
Nse55nMQvTice6HzA1qxrZfT171ta12RFeu9DHHBoWb13Cku8yMbMDoPBP2tl3zW9hFl3zbEvIM2
GLesUmiryi54jC9wYMvm+4fm1KIK4M8i61MQt19naa9FKR4yXPz4xdfDvxiC78l28iObO6Pno3DM
8wUG64XYyYuZsopsZ588LU+AjbxN2269RK2c8YSbkl6FS/N0mGo9yRR/HrS3ZxI5MWWiph9EO3lk
QjrgANWR2kKB0boI7p+ddJob//ofajF2Kw1cdQr18uLCmgMfcfuvR07w72WCj+6SRvUs9MZYYQzl
OHOJzDgcoG1DJ+f9++qB00I4VVKFBH1J6KRllmfYctpQXHy+ukpLEI5WZtwfvuPW+Xff5m/LLv9e
5I9lE97dBziXYPwme0VJY9q0POOIonO+UwR0qUl1sA0TRA3Sspj2Nd3UHis8WlwwSH9C/s2thH0o
3JTYAJ8shPAUnvmSkutzPw06ALh0UJmxh7r7EiO3gOR1sdKzy/LFcrbUvmS5SjeMuvaBDKkvXCRO
ciHKFc7rsCm3N6h7BRE/OPzTCUT8Uos9PpQBqKEnYe6jYa5iH/ydS5ECYabM3qav9KQ6m5tfmxBA
PZQ5S2HpWUKpj/RJH9OjS8EBNLqsHCGMDWMQSPUmidqxl9RwOY08FQR9XiDi1tEBX4eETh4+32OM
irEmTSiwzVkCHaJhP47oAzkj8T2SsSfBpr5oKferScfNLprrQrSxqlMnrwimE7A5d0vGWwBLZex1
lEv8itLi8uCsA4ixlBV7Z5siDGBI0u/q3J8ZFZuTnXD42EZTjOK578oyCRIzdmVLI+A5cCYVbaC5
O201ta6DF+ViteSpRyU3srU2MqzAkq8tOmz7x59PqX+LwLnfQTnQsU4ADLvdYdhrnXzhM1A8jyKJ
aND4PwS1hMFRzEFhOe/yvR6kpwX7tyVB7+Xtn6+sjg4bxeL13XeZGPNWl7vXQW4z8VTeQm+Gg2T2
eSaJHIe5p8kyORrUrq6Tdl+Sgy8k5SMBucsahFqMFkS1H3cBtnZkV1txg83tN6r7UUOxWz+ITxlz
FodoI8qijCBl0q8LSKOy6/W0QW306e0vJUK5eY8DPHBht2GTcMuegmWRKXoSbtv8+JSf2vHjlgqE
msQgESXA0Eom7Uz+gA+WDKLHuweepjhBJvOReK5seuElYzfiiLVd+3b97wyD3ub+gvGSdXVKPQwR
l78pYO2XT9RU88eCt+6Y4lP7ovsJo+Zd9lZNggDNCae9lIPL0poBT3CHNE17Kb7/tFTasCr2fkes
Gzyy8t4ohlMKkf4tso5GHTGqfQRa3bQOBytmvJBwQS2C/3I+s2IGMX3krQRskTbU4sj43V6NXOG5
9VG2ktV73iZlWzxzLsh9dHGrnL5g5MMb+7gsfjXXHHNRffENDUnlLuqQORchRoau+1FmkXG2N5/q
aPAddZHA8J1g4EE4XxJyEUbs+SGX808biw/YK6wjYpUA62+dYgEW+tRga+GUdMXX3ysRBibh6Zoh
NCdx11UHWzIsE20nEgMnQjBaKPtO+xQuxbMCsRgapfgUCfqBXieBdqhzWxOx5h2vzKMec4W/u3Dx
C+mLz172hYN7PhS/UvTLrrj5QkC4nfYxXsP7d2RYzG6XO6BkLp5ifdpdz0NuouQjTGKmWZO5rDbU
6Zg64ZgBi7B+T59TYN700U4b/15r2OkHP+YVCDdwZ0RLWi78pdXDHMLqJWCQct5rXkEY8UaGmtex
jE4XUP9Y4Z8V4hwCX5MZvyoD/2xJ8vNTPru2k4h5Sk5QkBa7qYGqAOp7Qoay1W/i5JMWDtIrh8o4
oSj6niNXItRtLcBSyfiIe4IH2r0lnqspUxqCxAoztOP7Tx9vLhvEBSdsBQJBsLcQNU97lfZES6T9
7dgzsF9lKkp4T+HiNzbLoD3n/OmmCO645M8GEfSV8Duxuw1940vekY/+7kMpkiZWQK9zaZD0b9Vt
R6u4llTlMd6EDMsqLNXTUiqzwxtNQut3cGohzrlp5W2HROTnl36XrDtfTAqmwE0/m7KsFJkffqkH
lJN0mHz5/8uE/as3z3X96skJKu+x23PBO6wkfZNj3EiSR7a4m1Z3w9wSsHNq/9yUUiKylnw5e1EL
TWDXkPKkQYmjXV0LOVHh3GOFmJMfA2Aol3/VBPsEdAQ4oD0p06fOr/e8GpE1gc21mr5PfhLd9r5d
xtMes6vXes5iA87lyKZLvPSeyH9en6W8O3ZaDGK/5rTtE0ewthjfez32EATU9w+sWZ+yFWMIRZjo
bIvLP8ZSZm85Vd4wsNhzHge2QytMBXHskrBjm9VklA+3yhs3AfmiEjzIXG9/MFEkjh3zTfCV4RL4
1LSS4GOuIOXla44BKx3/pLqmpZt+DE8ymDWqZGGRKY8iJd44yYK/graP9IFD33LnbiuBnLfxrQkN
bToWU5lFC5xBJ1uVBSGUcVqmb30KPG6WM2yDTDbLcKMCYzxtR3pDg94AFMf4oESwe6ryK0cUJu8K
RhtZ4qo6ckrCIKhBaMZy9Cyh8U1Nm6rJEJ8iHVc84aPVsOGOd5tK4iO94VQwP3u+nwod/r+d+ywU
c1D2roWtZrjJFm74RBn/1Fl4ffOKFGtgCTReZ8m6JAUKrMAwvOVmfhPvaxz31YQ7BlJdvBF8H/R/
i8c57SwFdo14KsryvN8tAEJvWTqDS1FKBU/HJVhjt0vON6HZn2Bvb/OYXd2kZpdN7nkVLUtPw5Ux
XrCBGG8GJVQr65+1bbR1RaDPG9ED0vjRtw4DCcLPG8lbtcyf2My0/Ru9UDXkWjXS8H/3dTX4em6A
5diRcgTyx2XmWzWv2eEOUf5MyyL+nhEVf69nMN3p1Z/h9hrPfH2DqL2t2IL8KHeuhi9L0CuA+rvH
SnxrDBW+4VGJwLJUapksyyYrYe3ECbgtSHNh5GMeKelGNBJntxqk17SEtUUO2FHl000C5W3jQ2Im
RhaxBrTFeOItffJy50+ATTKF3LBrh145p24gi8Dm2HBm/XaMynuLZPwQD+OPnOIi2RARknqMXnJt
tApT8AnHnUqYD95VwMyD/k41x5evVdcOKy+1DlpRWHJUVbnWSkIO0n/eWl64dkNE6zF9pWcluEdj
c2bWzmSTEYSOVd2C0p3DjiSOqNmPRjhKflMCtdKe6oVfjuMn4joGIV6aAKhnKbvqm5q0buHXp7aE
SiXvBTF5Qj7BjrCtfnPUq6rmeg/eg5VSvkGWdY8yHrnQEDkdtHqZhj5jVHDgUfksRPR1ok+kTl8a
U20uw7khzx2on6eADyMq/iSUJkVejUwi1CmN60pfJNDxaeDxvhj5w00RH8+QVpxed2yPr0zbCHk7
P90xXgHfFjmgU677druxWcrtBkU+ML7AVSj8qw5W5Qf1soLkTkAnFTt0LMr5sMczzDK0Ftm6yE/Y
9UUxlomiUdWl/FF7vNKoR6suceYzZG/wXsPbsQu2K0rm9yFxGurr7kbpSt+xlATZToAVMbEv+/jS
DQbj7tGhVKhPq9GegtDdHgftRI5ouBz3MuULehuV5xwdV0hbuKYd/7uO9f/xUa+ahpENwJDFkMjx
rr9QAJLFJzcP71XCGbuGbyieAGseCtggD5CSnYAIF2imttihTDFH9nm4yCWMc7c56ph3HiLp97YK
SjQ5KNer/KYyx8GNwsWoKiYMiKJsZOJnrQ/oZ4tQAGnTgO1fU6QOZwt9GJcuuOzAMDLxVWOAE4gY
yJi/SAZggg6dUCcYQFRrvNSAQtdgQAO2vQiMpBLWnlieX6WHBnRZoxVkdKgLJru2C5MIioBGfJAd
4amaauf2AAtJjdjk7HeWdw8Nz+1pB/C+67SUfsNxYP3aQPMF2/bQCnD0nP8UmAkLAtSRDA0sBhQz
D6tqjw1+6SXuJmw8rd7vdl2BaGQt0W6vtvUyGk0V+69oCuKnzyJ2x2FFiNE8KEWd2wghJ8+u13Yn
JNqy4YDHeKp71y63WO8b2igfsWJR/uP1S34rAiRkrruZKdPq6GGamKeoZp22Y5Bkk1SGQCE7b8gU
95p5jXEHn6wGUi+xIEmghn2zkcsVM5q8qHu427/oWJ38gu+dElgHw++/9fJP2GHSWnr0keZtAQHx
vCmsuG1OeEOEPtzEH+KDYtgkskzsmrVU/2PGnu1ZOB9/U0heDwhs4cvQyiNja+fgtpoEmhLvSQbx
dK8mT/sZmwas6DjtSaxcqoa2+nPe0Y4tNJrlMpKHymGImXVgyKctDByIJSiV6+mpkUcGb0cem91b
rdflMJbLp2cJUaP9wOOHQ4LyRCxlFrdSNxuj/vVmYI7G+jW2fVd4AkMWYzc+bfGCk+EuXnQKi09d
EHh9HF0CJBx9a6Vu6zekRe0wxTVDu4jFmBeJSO/7J0e7s8ERPX+HkkRoQiUGMYXiJkOWzUvSNGCG
uLpG0SQRwqEjWpBXj8gC69UqhcXyw2giJetR8d0KQ+mWeXJsy47+RhRB7R8TlnIg2j7s4ewYH06F
7XJOYGF/4sGaisrQNePpA1rpsaYHW8pgruufp0NOHSmrB0CLsE6ltwC/VnS9dwclGtHcCeU4C+6f
7g3DouI56uPJWYMzwrUh/eZo+LrfhXwnukEdZ2f5gc+yBTy+OQHi6U2AAqw/NGiOlsOqOpfhlLR2
0Tkaw0rzFKxMoR7GgTiiq9JNrnyvJJIFxs8amCA7fOxv/d8IkSVbQjWtn1q3k7yqYKYKI8X6M9Wb
hOKaK9EcJzauwp3jLuvJIybMjlZWIPriyYbgPmSVtxBZzXYUAJMo4DnWkJjqygYPvOLt4v3fK/2W
qCxiJLV2pivthnRsGr478bDAXFsO40q4w+c+TmAYvkGXQyh/izwW4UMbaNvG3cgbnGZnKV5mhjXX
9lUOcNO3q41mQSKpcLnUpLtGJP6TM/uVUHEq7JyqJkq449G75UDUAN3geoDT0aINJloRlIbxMRAs
LXWMSpy7e9wiQY+4YUY+Rlp9KWxsToSum3QYLIiy13rNh9wkqFYRMfIfgL0Vfq94B5b+WnRjIs7Q
zScFag+h9xS68o/lTZvoPzRxumb2kl2Bc8dIgRHbb/ZhJJ0XqubJsTq5l98+MqGusCRwrf6sTPFH
/vuZ87i8kr2RtxGXr6JD7KJ4KAODSnEAuyuhvytn8RQQsPAiQAt4puLPVAAYLC042tsmDNfvQla2
cnYUKUUzHLZYFHzqLIh3X0G3Zd1zyW1gpwRwWrjszoDgDkR0TNXuFD4VNppK/Jqj4bDLv141DaPo
OQSEKjME6o1qGZK6z8n6UvPPaysi6BOJklunVAdRLgGUBF05BTf5CeHa7/b2mfJlsq9YjsmOg+rM
AE9Jfy6G3zQDsEG2n5HPYDAuHuT/G8YYXeSA258wQmdEXmukzrx0W3ucnVK/XuPoinu9r/EUSt9K
FsJDUrjoKXHDFVtLzZVJtejVSolhj0aZN82/oVTpvnc27NwIrPNNpQRjUk5frzz68IvxbQBRxbjE
WR3r6kWuM+u+tnN9MGkDhu68QS2qZPvgXMdf+Cmcej09/wznOdhys2rAqM/5M8HmvYVzaS9cpMf5
pF8GJnEh2joQFQMMZ9DOM/GY6iSrypuj+Wlhru82y/vMT3SXevSHGwC8+76iSbRCVt9JK6dHNINx
pbsHh1HnAfE241bEUjuzqbUCjlzBZYh8tFt4mR2PfFBtYhs+5wF4FGHApWUMHSHnqSBZOWqCxw7Q
iP7hIgEqt5QtN8pQ01srwK/Htcs86Oydt2iZCEoc+zv2Pp36S7Z13Ago8phVmko3D+rpliT0PoZu
27GmJEKMUPRJiidPIoRl171ZRryRFVs0i72JXBDdqTjeZIn1hA6h3fFsrvgIe7KawmQbXI97skcQ
J44qjNAYRj6CXF5uj7l5CyFuPUBNlOJNDj3exb4f4sNC6uxcHnO6Z3v3NWegF21kBHaexrcIlzn4
MoawOHmW42YDykWf5ry5rxJwezhOPhbQFAe2TfoImI30KcEjcNPhPHYq23BpXbtX95rLlfhXOGcn
QP54CsQd7wokmtUSTuddaEPKTaH6LH0EvMpq19q6ZUDaeqlUChdpjJjCUPJLqnjKUPP3K6q0UAck
DpN4at5rdujzUIW1KIq2caznzz2jAUD5qxoFy63z37QW7xWqWu0eVXlIkdj07RAzlZOtOUyhWlSl
BQh7u2c7y46qjNdzdLIcxIds0sEbFcegifAzYkti6KVvxsqrlHQ8UKhHboX7Nc7wUochOQuASRIF
DyGyEKjMFa+jAO3zoRU6nXGyFEVICvzmxHd2swZaHo452r3Z1x6QA+EJNBrgWu/WAbCU8E3F4xxM
8zUpYVJ8zO8IB8HPo3XfT5pCF0KUPTp83Nfe+i597QojP77xhO3UdHLlCbpQdSXxa4VXZfcnJLGA
e40XbgY0e89+4o8Yz/Co2K4epgpxEbNzYBMawjEK/dEgYK1cEzKwXrlSWapEjwjhjDLj3sQTrslD
K0TIJFDgV1q6eIhTTpZLzs5WIIe2n7emDCyT0MtVkJG1uSK1Xz3I+In3A3OsQtnC6cshOl/4yUjW
qUbUF2iy6KApN0c9BIKPE/TUArmGAR+WUKAdJWdatkmGR69okBn/fFxwQFiEpXY1YlhJ1tXvMYXr
S6RCDg4kodhObaJ5hU8SM/FtvOpf3E/iWCi4G4J/Srfp9fNTOlV3YuTklLlxBGFZyhVfEW5j9/0c
gkaDSvWgr8LljaP/f1lJxT0h0OFMrH2YTu7mF6OistDJ8mAHejo0GQwVvDxzRMbfbj6cxvs+0hGf
vMjhgwTgnK1ZOyqydBqcytZoCrFUacp0gtVtBkFiwDYgxtCDAsIT+iL5bhfT3GcJDxMcaBeqwdhW
xbDSk2/1ZqhcnFTaWTLg1pE9Ur9dTMKbH+XypGxLcGzpPaTkDtUaQiW8Seh6s1/3NxutrCBxgg7N
7EHuwCqPaYbThNI12C4o63Rq+8ieGym88qui6suViWKvePy3mflvukU2JYn25yGuO0U2b+QWe5Sc
EzqErLvrkhA8EGkq91FIl6qZ/KFz3niipLSnTH4427lGUQaUs+aPDX8xwJeKfWuEMsFTI1myC62S
ARbEbo77Z17A+FRM1TptjCOLNNgnbMWLoL68XXQP/cdEqDlGjkTZVdSwMCHi8ZbRSX+53Q4lM+gf
U5MilDtKeb2VwjXnIzNlQlTfIxWDyuauqi9sEEd9pXBjrCrLhguafxHGSQuoVZ1GSPdtRMnPQoMU
1U8lfIF7mYV5xXU2ulQeChPCXEblhwSvb9hgYqi2jkbIEr9gQaJH0pncHzmCtqgohFFxWr/fqMPG
hm4nzGB95bSiFm9riCoQ9PVooYp9lwXEbiae+vZEJWxb3yo+UCc5sqLBkkSYrgrtclpAHWrb3h5u
4H8pl7PYlb6yo0aG7abatUQBMXWVM5AhpmM8e78OrNc80u142Koi6ODAg9qG6AsCYaNRwHgXjQ2g
OyBWXFdLVtHs5yfmxT3ZvtkHxub39BszFe3lUGxNLn4R8hr9aAoUnM4k3XRURsoBRNRp1T/0D0Rn
o+6Rx2Ik4FaQ8TFvqoyY9mukn1nwBzW9jgnPYmvFcbaYlTmlM8AsTPs4mBFJGWi0XkpHy3eCnnmf
Kvfo1uG9GR7uTV4PgX/6k3eG1hJTi8PDSaccsQrPSOWU4Xa5PMg+xwPwP103geNa4eczA6auFg8z
PXVSVA1BNcH+or0P/QBjlWIFhWIRcf0EG2qfxkSHLNeLBjWdTuILgm4qFU3zpLrmdaoLLx8K+ol7
owv2f/UXbXN4ly6BYa4ZLGSqLvTWfv5HpCTtaHmECIGoB028GvkHMadT42u7MCBBqsYKQD2gUPHp
VVMy7YbyGsnXkpi0MgZQCnZViByoysbYWUOpUfntqM4R+F6fbKd+1P9fPrH2I15s5e3kG6Sqwyda
R15+3ZlVA67AWbL99Gw9bNGny4y/wCs2ZqL5bG2Ux9/70TLqXPVBTB8jepGkL0d1RN9qPmafGyvG
hYFBnzYzmYGLE565b07BKGpkbHoH9vFnwWP2YLU9+On570q7ugLZNVaD0sW4/HIXbSGjvA+0Ndxz
eZyJm27ZPgFsWkkm4rVkvyJgvujLCCVAFJ3oVB+wc0dSTSeWS2ddc1MfoS9863rHY++Y+CGnftaE
G0yUe9JX4pHOkImgRTdF0iN3bINGG8MBOL5wk4L6hw/LYoauZRbmgVOVsw2/sQqink7X9DTBOu7r
SAA6i+Ca04j1QMpdF8GAMkOzJ33UXHBlXajrSLYtlvQnHyiKrWUgc+dKOI+MgfFLXnUATNbBd6cw
1OCSE814tC7AWrdaICA9JEbPBQ3LLA7X6Fn3uiMDvB63TZSWeDL1j/hygyYYDAPze1HU7acKVpZJ
/YcSWzNVMH6pBOJwIJckO/1cxcidJixcDbBWaKPiHfBCpKzRAUO1wwzA/p0pumY4rvedyZ4Uh71S
Uy/qKALyYQNWNgRjkOPqyJACGNQHFUALhfmQVbGo0kRY0mHlIMLt8nl44DCvv6jNXQNjx4ySpzga
rWlZo3/TUEKQI29B/yngTvR/AZC/QOtJIzHwMaMNN6ox/H4AvqG6I0Xq3CiyE/fvQEedWluFgFJt
zFbcgu6/M/AFzuwmB1RMv6Fet2+GBRNaA3VAQ1M9Phwd1qTMDUSOHGk3Hq0yYyHIBC7bHXm/xtTp
C7+LO6NU3TiCwLVIf4aNdvzMLSe+n26mAVSnk6pB4g7IzAeeNRkKlEhryAHQBP/m7QEw2ic8a2d5
siUus7dzUHzPLmYDXAQ2EsTdipci/TZ1zaxT2onOs3DJsxZoPuH//MiGfpjKgql5pSJ70CrRMUVb
jU/6Xr/FmwNBXhgOtNg4DRLceNwek9Z6yBSnSAIz/prIww5o6FfeD0u8sMvv6yG5IRuK9w+Au/e8
zNyfHg6fMFzrk0Mxn9Xn4aETlUssIfkMybmstTF6I6qOdrY4M0dthpo+wwDnoMkY+Qafjs+M8rfz
vHQg8+8CgLoyQ+THV5JNIsjITbzWylXrKfNJnmQ7XFf8iyBt3GQnoNLKc/rJtfcGHvClP9ukWjZA
CmsiNjiKaJQ+3imiE6uAZP29VZmgYRdYuQ7iKK/dvhVNtluQrJUR6B+gONeOlsiIHMhx6mNHN7E6
9ZrOt6boModMHy9JovLYg9P7gDlX1lihulcfEIOOKFK91hV26QGeUCucND7C5Mu3YsY0+H5ttXJk
twkP4XWQjVJJ4wIL/QZY2tGLcBryhvxEljKYB4NhUaiqNGHSMNBpFKl9ZRxcYCdqrsflVJD/dpyZ
BTaGDfTEEV1S1dzKv8t8aGjJ/3E3vFqgEXmVcVdAKq3hz0wOAuA0rAWGNXfRveJKKb6brz5R1yph
2HMrYAteSaYgEXEoGO0Xfthwn0bKKjXKw5zgt9yP6CNYY7hxUfLQ+GdUkoRLvuck+0AKQ2wtm0g7
9iRCc52mYm6QWI2dk6gjKN4rwgytksjlvUuKno2UkiBqsZqOqW9piPWLkVD5pNDkaDlkZSWTV6Xd
CoUtXze+uNOjt21XIPLexUhoI6Brvgu9he+EoSuGD50LlmHOZ8IOuy1xzuTWN+VEbIzDbo45fcSu
ltkdMK3g1BHR+vpntPyUn2XS3Ji2ZvmTVKtFTtYFUXJzIbFPevHxn9SbFfrK2bAS97ASsIFlyHpW
7APj3/37k2QZXqB57paZHQ6XjHkdsbnYU6MHvMdkIUZh1TpFk9+HTHb7r7UjxK3lG+DR9ZaXv/i4
FDhGAmZ2lg91sSOw4IbtVbr3RGt8hgsLKOJRXo/OHKJW+3W3pMeEFU89Kq/X/bvL4CtLcnBoqs3C
gUihBNBs9LpMk6BFRj/K/Ia+aRVGjek5kvki2slzw3pX0c/U9Sfbk9pr6GC/8EQWZJtmdzuuoMjf
6BSWXhHppcExV4AEPPQw0K7h/bJdffDTrjf7b+fdnTIQTdvgmEmzfUfueIE8xNVJZP2165npgfoD
R5h9sLpTcia21xVMZhfgEFkvf16rMxwguk3WH0Y1j9VmZVcThkgz0cEtXQ5mXSywMlAhsEK76a2A
DnSbF7H0nWqFFOjimQ5EC8j+M7XDNqNAfxy8QKbXFgZ7c8++pHRDHIo7qqU+4EitNkDgzQ0bVt0k
y7jbOZObmJ5t0JGo/oBeZoHvwFQkaYI9Lnn38BR+RaTrkGuXGCHjI/h9btbISyToeC+y6qawL0Sa
cbVntd5wFUSDcOsaGe7L70kYD2bsEW7XkGxuYdBSuAfADYs1AzpJram2N8xgaGHOZgM4R1A8bc3p
/miA8aWFh+8VS0fl7mEogkuY0/1g3G7HdgG0UNK8Cw5IuZe38EbXFWaX9HpM5TSj1SR10m31omx9
8torkB+1Y+I1M1MLthfToxBX275G/fW5h7bTXMberAa6vA6Q6Flszn3s4krfTqUXaQ5wyLR25dTa
PxfApFiaReDZABfGnX8+Lq9GMw4D6ZeRGEpUkSo5Tm+bM1dxX/czlhshZ/or5kehYrdFgHaX8EMK
X5RueSCuA/pw4BfiLYphvz7HcZGvi8PrL8Ck54Az2CnERdtIXiONhZK9zJjZYUbVkR7uHyBnCcpw
Ld7QzHl4K4w3ewqtSkd8oCA+mcGr/R7uHy1YQ85BmUk8b3NdKBzLSCSAkJ75ONnuJKwByxwxTOr1
OWPN+Ywbq/lyMdMDdCKuVkoihXKRJeR3YBt6pEH+XQ26Vdj24lB/s2I4+EDa0ZQSGkLJRQnQOrur
pkZ39CE92MH/vmvFE1DIh1j6Xj1hJAP+sPSsnFcQo+pxWRLhK1ducIhgglJJPvAnqLgWiUJZ8lxt
gUOQrEldxwwc/vZQjadjICkCcqSudSgEQOJII94IR1bz+9nTyT80Btxh8/Z1v/U1RXabbWcYx8E8
01D5v2qKX6gUrnIQlVGpINTD07rgjhNxI8ubm7FFLmmEOcYV7XWUR4PMT7NOG6kBtTjj7gruQ45m
R77j3CWDUHihh3gUcHLq04UQVlSHqVZiJuG1eqLm5N4a/uHSTtv7zqYFQBppScdQUoSa4Kzobgk2
C3b6RTPYw/VTEyPZhXyw5JfUOWLYbJFvg+k0R9PutPjs7q1WyVdhGWjyfwN7OExwcMUt7kqjsFX5
/FRdMC/6baqF/iNeOj9M1HdQQw/8Vb0TYxiqYz/ovMMRJsL4TmNksplH+6UlqmyN4BAb0XhkGT8p
PNFiJiuWXNjcE+UY5y2cBHxLNrTYqlZh4/NUchCbJ3do5tjpB90Kk4Ppx1Uv+bgRz3KprNVn42ZO
6b81e9EBNJSJ8NyneifH2aJX8RrLV+v3XtIWGnradkDftR4l8i0ivsp+jUY0ep4XMi/KtFeJIsNA
+5WE025rcOgwkF8nF0FNkVGz5ZCjz2LC5M9dVK7/2lhBqp5CxQIkdafkC7RWTmHXAVxnZuWVCelD
SOjqtWZ0n3KVk/D05Q58Pc9Sj4wQHMvxhBRWkbsUHOeMHWx0U26kPGbejxwSOJgzbyK/PnvLP1mR
ku2qfQHeKOAvZaHfrf71hK9XTTgG3dB6jzrenUu/8Lo04SB4wztI1g9clZQz9FCJnmb/Tg9XTiz/
EkKwi+C5aR9wde9vU0KWv0QQjLfBvOEQ+UWFlybR1cIjbCvEfhoFodzeDzVvHDyci3wVNiNQfA9L
XDP7tH0vtfqoO3VsINobT901zLXG05L4QedraiDMv6sRdPm3GZsZSsxMNQZ1qNIEp/njvkyG+4ZM
ghDugGGnex3M6tMy55PhhJ1J6rTDOZ+9/KkZ14rKKgdcHX/ewgVIRa+VFT1JGEJlZMDoitwy7Z82
qhBQOLzmHXeszP4L7In4+QNvj6mRaXpI785KRtjpSTgJhu9srAVZzeYm4YKUjS9ecTgtHdHwlA80
3L8980zLHReSahhYrrpgSwJp220IhxFro/M2ingwQAIapGnSN3yTF+/Z74GLiA1ju+Eu+LHe1i3J
hpElwlHI8DGYiKm3/EqnxDxFDIuqKDohk8RH+/+kQNWaFsKykB2EPWAYqPpnMJXy1LhkHQAOcDDr
/3s/2OuHSHt7IvtNOI1JjRrCuBh375n6CddN+kDzzjidn06czhEGMQ/bCeLSRr7JLJsgpaPTLVBL
NCTZIIou7VrWyYFogOqc3jNooF3POKOXx+BAGHpskCnkrQvUplqy6vKwejiLNze3QdYi5aLUEW0K
u6Gigwabzf8PVwvI+sPQrt9F9mC1oqXBrGGUOmuUnH2IWaD6de0guJ0dZI9j0l4mN/wj9kVP6+jD
v8Wj7gPXlMs7tJ+v0x9ZtHqXN/AYfC8biv4Iuvl6ffby8XpmdvrWw2kYliR7hLOxDYX6rs6K+DQt
U4LZeEni9Hf98Hq96l+JnwNG2oY7ZXKpRpznI3CBVJp0oJKFdKB69LSF3O0sh1BAuOYGM+ZH50dW
Uyfkf88GszmICggqV/zemmr4p1afxK8FpRa3kqjJomR+puxP7jslLWPODii9dIECifQKSa7NlAMz
V5oGeYfgrzOjTdYxhaNlJdkYYl7Pa0tOVATIaH19RILZwiAbJqEV3swZS3937/39DWkDUMQNEjdQ
U6lXdJHHADHKUCf8INJX3M2fLLLmz/oMK+oULsdQZof/NBtuRFG7nMIAFH2WOknIkNKvvBNk4Gid
fKGawNBOx4HLLRyQMoB+4RghOtkW1i+oOp3kW/eJra3nW1GyEoa31wfTOzYAA+bllMIrh+DjZFjZ
yY1A6NkOIiVILoX6dX97wxi7OOUNoykWY7bE9nz0EcXX8Unn7JDY3uYHo4tDzt+jchz7rN6KWHVu
GSV6EgvwARdyXfBfXnusSJBZNqELqv0ViNyMwHHevC6l/DqFIYv+JaMGpksu2vOhLHa8hwmdyfDN
UH+by46O/lgzbYnFJbOqnS/kgiF1R903kcUqgnPotfUaUp3jHUxIKoBrlGEjOKoFao/h5CktlJCq
WrXhPrV8epYpfMUQQLycVxu5iMxiOe8GqJoOGrnlou9wIBoAv/NApgvyTwSycLTJRi38Zcr7VNi/
0KK1o/TP7g5kzbUYNJidP8/fSAn2TtKNwdD8Y1rkwYlmirAQ4rUC22LwOcSvQXSVfdrh6PnvVm+2
q+x0Q2pQ5J/HAZKhwqCa5xZQNWuQWzffWU+48lju5FL0cKuma5b+MClX6m3nQoxzGxO9mQmbdRVl
CBjnpqG2P81rL14dN9ALtWHoYBkQi7xQ1p1kH8N6Fg1aMJiEPrmf1K9gvCxLexBW4SU/w82/uAq+
3xOm2y32+rABM0xOSEr3/hwMRT5vo6PT5Ynh4aJ/jfizMgRqui6KqrawgBiWsTr7ZmRK3uTvSV8C
6/S5dRmw2hIZ1nfNkBVDUA8gk59PHaKvOeH7TnglG313KTZzWGPSzfISjWd6eF720E9vQV6H7F2l
pLETxVysDQBJ8GYwVRtJbpQqCsL1lQsG9jADIPXqYC5l5Otr30J0DIteHcK8iokqyzeEG6u+ayD5
juZV+kqAl22HHEbXpAy91CjquO7ZmCeeBL5Ozmj25Gw9EQEZXnZRxFCWtqZ3ZG1E2qsPmo8YeoW2
t0EblUjHQabmYhw2yOSt8R6ICMqJxFuVxHWmXpVIbUQMztSbc27NsmnEPey0aCy3EkJjFGXUa+Zg
OrE4o9wirclbXian22pjFLZEJczZlY2P0lUcKB+utO3zzL8Ty7DVBPT9P2PJZ65SFFjwfh7oOhl8
nO4UHjNio1Islo22QB5AzdEQFvE50+4v68j0DbZ4lLPVjDzBbXkIlfQUTwowOoVLqjCiGFUEpNy0
1P6eu4Rc+q+qOQnd17dKX2Tz2tefK+N9BpDaFk2pb8HhSeNGnzCxiRpzPObmiMgp+PpqqxDX6afi
KIbE3aEDAIkHRE4lXXmQkdnJquxaYE0gd1KHjWNr+8R0KfejQuHOqwefutkj5PC30Xx7mGyO+EPU
8sQiKAtRpU17LOgVrJpZHqK9o2z792k2yqrkH/z7VvwPa+yqOJ9TPWGTTk8Ztn7GbgZdLT2kVgQ5
FqQ3AyGGb7tiNh6vemHPxjtEWUsSZ2tGQ3H+YtuO5ZmOjq75Xr8p/nlPiBM0Rf5DXmxUISDvKRsj
Spf2+SzqpxL11AuI28N2vJldK0A9eizf3XKQYGEZKHL9fnfBHSetkdspsjIbPzb8snKKKA3WrGYz
jZTb5dmfFPFi/bLPqmiMCy5RHnKXiOqJAdvRyLaJ/F2d2I15jJ1EPhjOWaayh2rOuWDL/azABCEi
qr/Ty32gOtQD8FIcupVvro8NWBzFT7q7qxFbxTMxRw0LqcYWyl25kDEPx0NBr/My+pzXdk4m0QFg
9Q2kKFK24KtyB+Nt1khcGs+BQD92sMiD/ZIL0gCjAceh9FGnWdWQSUqOuIj7ERjUW05b4Xh3+N0L
vmiNEEEN/w/PsBYYLiw2C04ErHdq2vox6k3AQMaTAAk8T0MY4Qmbj02zCk/DRkiy8MuLe+Z2N4fL
mK1AXtZGwMfp1zRnjHBWSRQBjjObv2Jiq7oel4akDtDYcjlIkPRyOiT/aBkfnL9FLyn237Nh+g+x
n9mLt2Y+GkYkIx/V9uYqjYIelxjtE9YhNUHR+BjkOgjMltcTpqSZQFuoJh8EpNFAA7ySM4QUtKxB
is8u9AIkv+BHYeE4aUd6L7+Mb/dHchekTqX4Cy9WfQW7xGmMRueC9KYA1QOs4e3ob48LxCU3bKuF
cl+zFinVSvROIsqyUGyInnOJcULF6Yoe2DUK7679c+TZC6e3cpWX46lCwQ0etffXvi0siBykOV9c
APOfWMsQe/P/cyRupeln7qKnShuy0L/YIIZsHlJFbymGt8u33fQPSFPoH2zIXR3Yk9FZ7+UxN9vv
1nlouUMJ/IGxwQ7N30bJSUfjNkLQ4TE4SDahKdglHmH5LHTfJCUEej7jucvMkh1T15GJ2VRUlasj
As7PfYoVxrkvgs4eGQ+JM2BS1VNnsyBqiJ/LDkjwdrTFv+x6YrIQLaU03knS1gA2wm4gqcnab2DD
I4gkoTNJB7kvhu22o+Ifio6QzXcys/1FnZYj8m+ZFpPkSrrvPseiTvx/8rEKfEX99vJnDD+Tlsfs
HfF/M05zogVXGdV/fJaTDhUE6ycRi7S1XKE3VqOZ5JylwQN0g+XjUZOrNtw5SMTaBkz86AkhH6+y
R7+cHkfPD42WbEAAV8LWGWpPpRtobaKHA+rIq+FrPLdht1VlEXlceGxnuoWhS5LD8MvUSFqImF8u
pRRefDyBXwNym0EDQB0G4Z/M/cOqFYVhu/8zCv/DVVgIKDDs7Ahls6cW1xja+k5ziRhOgXM51wym
MlmEy0nRM+peuyxPdV2Eu41o5TeeQ7OWWWO/w2S7RzGd2tg/nRJPWlCFFoBDwwDdtJff2bYnTp2C
tb0MbwCJxkY38EkdIxG5g/YkL8gynEdcz31yKfnTpwe2KenIQL2ZAPyvx95gsPmNxnUY8qOAOlxL
Cwqr/iZzaY+nNuQl4N2ynS5BjuH0cx9xznqPpsVlBJ306L7Awatk4wkjCsXa2edmj60DMt47qfNI
jQA56Vv4DtIIhN4gqteEm5b/xmGFiAr5ytMJ7Vx2xsfysk8V8FgKdOjLmO2D5rcR8wqfkI53zUcY
1pGbEj6MCsakcERL6H2FQ4SiwwxSjzACw7ADWeAuULYhya1jMbB+2lD0FldYS8/DliM0U7yaPVeu
yAG6/0aZUgA7sGkZwi2XuzVW35ZhsqG+CDwa1EFF87DorgKjrn0ye+tV2yMRz017Eo27LtOpEM9q
LwoV3aqZyLytgWegn12uf9JTk8jJTPbSaLWwOS7LQKc02MiGSXpwrmXAB0HfGu7G2dm3sbTMB0Ww
/vWA45vkEdUiIj0nr1MKXS4sQqdizVw3R3q+sz/o1yQjnbXlI8duoKh669cV0tzGGAaY0PRCjG3t
kM1clDjHJuIpXb+n4AwbxnyvYkox3GCPx4tNcBxGOWaBtR0wFR/NQ0gXoZniC2Gz6fQGhico9xQl
OlLWCcCOzkQpDPimU0n8VejhTDsrRRVCP3OTsNkG0U/h+WR6mSQuFUMCqfcWqLQMtg3xtI2nNXjk
LRmgt1tNja048bOvzhNd9w2w6e89+PbHDSZcwzLI/oD01BxifZSqSPBAOJAlDPFqJJS78lMylwov
r/TDUzDNFSUiha3unRFdRsJkfukyGWsOoinLnyCuJbx8gBkFHwahG5AWTbbzFP6Ia365HFORBdEd
EbycEPjTUjuxPEd0Zq4m0rOH5kH/hhHBYE63may/q1JLWLDr1CAk8duTTCY+s8WMAC3YR4zejPAz
13MvF+lAWeKGrEsQdOSJsZlXlaohDFmhtwtIEPJeTg9ML+R6AmJBoMu36FLwXh6IszDMfxqpyjEi
X6hNLvPxqtvtcs6VfEI1eqLaYVVKHYISraoJlFLkb5kX7dBLmbtedy72e4/PWZq++dHrm1Cn1+CR
tORITMpfe66iJqaapsJNqs/rRd4GODkzOEBsiALn0S76JQcsQK57v5rUKcQhfsIHnOZgq4bfgxz5
xovI1xfCelt2UKau9GVd3kta/luwTsYzAqg1Le6jMVqdXaSqAUx/I3NyAl+NNzBrkswdJdjgXPwt
jA4APr/di8Xjssaaw0S8Rdyz0dDuSO46XOLvKipe1uMTMaWUifr50MHonyH9JQ3Jdk5qADwMIedb
US/xA0iCvw94U94/1rdZngCo8tFdaJdrUF6zDvb1T2aXrpi6iXgTD9kJzUpU2VyKr1DzObRefipS
dN3of7eWd/dG0UYJMj5SE7YTdKipo090wO0KHWUBBy9DhqsltXTgmpxGf4Ob3+cSMC60ynVIJHrZ
kTJLi78C3b8+Tnf18Pu6KZE0grCi1mqf9E8bH6WoS6V+AEy/jlOi0D/6pV5mNW7gXk4hYHkGvLaC
z/dSgOQLMuyF01UcIYsQaCiqbZCIQmV4BVC/guErKNp8EzU9o1JYZ//WVxGBrLtErBVJoeCs0jB2
SaGHk51j2Yn+nRozkzix3S0oRZyDqy04MU8AVokeOEDxzpXtcBp0aEpVezFGcgWn4FvuZ8GyCvFd
UJ6S0qw8u/2f16cGYv2W4Yv49WpwEI8YJLv4XfIb+ces3G1Z1v4Qit0B9XOP5FtiPzCkzJtTktP/
K75wf9oelHKuHuYunDRgfB9TRFv4iO1Ke34soqOMpJgWCu9TieLOc2QmD8ahl+TYfscXHIP8fPZS
IrNxzOpj3/VqVJRnqzWdL9xM5+C7V5epNGEwj6fWNoH0jpMyQ3gV+8Shgxo/eNkGegd6fr9DbVJj
+iOjEjI33JoFMeViKWPHJdp8JPqcHMOAKBBhnP81eSPbdGI5N3WG0jH3DqLPpdiqQYFCwXHthvkC
3uVk4bjVL1i5UCVtRE05yPGrwzVeLjhFpD58plwBiqPvu0DE2MJ5UCiHnEFrwvCdvhIYQPAipzPc
syhQV1prXFJpwCskpWAE/6StLCwTf27V3G7LPHg6ZCH6/3VQLmH64q9HNPMCzg8OfItsbpPuUYjg
2B2gT1fZ2efn0iTXjWNYu72/SJ74MMNMrRLK96o0TAihTVeAKIhkpcRe7hKwF6obNOw/XyIii5jw
zkD1KAowFKPnjaLzIKS8I8LjpEK9hqm1rLL51BCmKW79xOvvxFFuwjm2QfTvBptdpYhztqQtEux8
1Wxob57FkHHSggcLJKp+VtcXD/wzyL5HLaR7AOPVqNOAGDujww0E258n9b8mTYbZ9A94ks3MXrlQ
X+EY8QLppu/hFFYEIWG+evKclSVReIcDlt3MrWJ6G37O6GWDYkI+IZKUhtgzX9HjkDlAh+mYJ7s0
SqLk5nnpsm1ZSAd9/GdKxHuH6oe2A3hhx4Fy9zZfJFkd20FoT/MLP42Idnkal2D29fn5PlmjKNkU
K+lThK7yqCe1newyp5APrvesZZtWVweWWAWnXGFUdw+x9SPiBmTcxRLbmxWh3tP3ijpSXNwysrnn
/TbzGwuj6Cgzd+iXWsK5SnXvX+7PZBcZXsG7ZH0g+ckEak2tV7MCaomu6DigNRrKDa8tkox+lBcJ
/45ykB03YzomsdJ8mnCCIABrHmt88i34mr3vnEHBBCAFMwKomeS0WG+TB5dQfXu/YWM6aR8qoVeh
Ko7W3r3uQJTsCLX/K168ROmc1iuHEZT8cF0eTbfzDB0oZBmWy7FT9tGMDLzQYnM3ed6zWGror26E
rw/xIapwXBAMp33w96za09mMiMVEXdUL3QSGd48n0eRlzPJMxdFeiMuGq4LOvMbpP1OEnk4pET34
ISJreMZcugtjMfUoPmhRIz/2+7wpZkGdGLn3pRK0UtersO4JWqqaPffjeJIxHt59tXRULgWhnyHk
eY/VZ3ixY4XCtJQH+5HmNrXn/fXh132WCldz6wfXVhSN3YETI/nnLYO4Jx2zT3Li7ACK3rjb+nQ7
psTswJPevis69ooRLnjzFa2U6VVL5hX3xLZa9lCyN7vvWACjyBCPXB6QwtouqPd9zPqrLXIuqjUW
9tlOi7uIcgokEc6mmAxVt+8whpnEFPPD/umBvZ1Qz5nheT6L2b/9XQSwsntVsU5+rsK65tSfR1mb
QhI4K3TytJVG/i5uTHq9X7+eF6Sh9V2Iu5p69bNuWrHFzFqgF7PZyMKgI4EJHhFkNAXcqcxFTAfG
WynzVxrZjhP8sGDLxIrmn3y7nP9iqBwDcLsXdW8DCCYFnI5D+xliAE3dSMsb73K1BY40vviXwfaW
JmnlkNb/Gbh/la2K7JDoPGXTAvV2GZzLOKbk1X1UxSjFZWfptDKBlZXCVW+jfsW92fs8OTtO7Olh
9IFhlZHpZOQlzC4Hl0ztLiKXnyoPJdDfSCiBJC8ge2XiS3Q2ddCVjsF0ZL75f6iYOk/tOfIFO7vk
afq2Jigp335FhOz1dBjYKoepJBkRMftvxfgi77Yu4gG1OgWJeqeDVfj5RptJ63gGl361Kl5D235D
6ZIDTFfeZQZJm908o9EqPv99gPdORbrYiuj8sojEyyT4m2gx3JaRdiQeISGeAE4XQVuaxZi2B2PY
epF3sJ+TPgk5dzHO1yJ+RcY1dn8Pfr5OcD0yICgI23GcagYRAgHMVEctrN3+jcD/Y3XheITE/3OO
FghfwrRbNImaIQwB9lknlDFcqaX+sZxWiJTPXyC+SKBK3HQYnDnFSlsJDPRtytcXXqm7jDbIOXCQ
6qO/zehqsGfzCZdo8CE4WzkB+ILxacjBQgRBbylwzgS8HVhOfbvffMTb9fnoyU2f3Vl6nCpnljHi
77OGZk/DJu87VR+O29M6RR1sm4rpWB5+2ZS/lckX/qjokEg/c9ydy3+vv7YadqwKneKk5xiD9X6A
xYZf2A7awsIyCtf2NgPcnO3cdZBx7vnGwbcDlkXcIZCcrEWt2VumagRE480ynV0/CYRn+2jFfYej
blVJF0Vtx4FW9S5YDgtCunkzkEzAHGxrBRi1T5KdXO1FvRPZviyuF3YXN1mXJOz8Zp8pblxoIE0G
aPjFOPXdsMy3WOT//eFoE4yXzbux3m6sYSa9qpAEEOVsmG1K4ndaNkepjXn3HhrUgEiudq14qsaL
QAd9dn3yigppoJ4/lEZQJ/sV2sknAHoStrwFltl3lZup4UWSbnKWdewruEUTS3kFduuXAm+V9/AI
IFCMgABnAaLapYhqtHrNN9g20Whdtg7EOJ3ecC7eqZM50JaJZCY0L6sNsQHMSa3mgYra3VhL7bBz
/7fKA8oq0MXb+4GjQYSCdqYMjvHtNS/kJXUuJYA42zHTHIISsrAd6y1lo5VH45ZSD7K2RZok06WC
YAkAcmFS/dIp1US5trsLUI8oawmQikT7jiwswXYUJD1vPnIWVo32d7gk9T4lK9KUfUWSD2IWZYCw
6k8St5NkkvE6UWu76YVqK0lOaYKEleUmPK7mcasvHpjwwPkOJ0FEy0T0gTf6KNiGoP9UD7x49dMA
SmGe181QkBgh68jiCFj3DqflvEEhSBnT9QDhk3m4DKkBntpX3dJzpP8JXgik0x1wvQWR81/mXESl
M3P9/n4Lhud/lX7UXw4l1Gn98Mdpy4K+GfrHoWBwh9K8fLr+c4MXgiAsdh8jxbb1mFFWYDtkPGNt
yAQnTKS4ucmJU7yvG0NZDrAlm1gIMeUZMCssWZ4k936bGfMS2zlxCWNufLTSPSVYkVkMzBnh9Oxt
ic+w2rr79C2JaA6ylp7utXpmwS8HRZmISfantcqjT3yqmA8g8DWVBNG5uh1kMNIFVf8Z0pb5u+jh
krR0t+MIqUwV5Gm4FJ0vOrYoMYSRxbR1sG+3kZXrIUPHLgmBgiRwtP2eM6n9/qM/kHA6XcpljUJg
M2ct971LFd1tRJL10tB9+jPDUkj2FX8mGuS47jDjbxzjayrZ4G+RI6/YEuiD3Fcx2NtIdAkM2HBF
MAG9YizwWgIg6Wp39DVyA/DKNZPi1IE/kvkDZiuUv8jplco4HM4XWqpnr7rqChNWWz+vlJiu4r7e
OzuZDy5k8ASO3NG6k+2zrIAHysLkq+RXJ8GjSXcxzyQt0K0FkBm0+6sDLVLNMc+cXvtEykpNzlnb
k56XpmKJg2Bb4Pdf5AOtwh39AuKvzhFkF46V260qff8zvIzGBUjoz6k6Ka3+TuciYEF3dK5r2pyS
Ie5nNFJehb8qkjseXOUDcigIcuX46zhhMPJtA8FghDdqWtfgIx65WT4M+6vch2z+fYdTpjm6fbba
92t7rLwDcWPtleAa3kfbqO/y0yYUrZgCVKs9QE9X8lFCIwD6oXwsIEwy9c2585PKUoGSw9ThgLct
Ilp6LVEV2Zv4lh0OpncfvLxzvCc7Hhg4ANkRzcIqssu31n3op9AZ/qlrZeNq0+vQ0OErju3s+dCV
i76dAOsfGEqkisEUjkn+R8T+t8IeYrzk9ktwRX24rv+XADKZl0Asr+EAo5RSiHBVPG2PwtvRafJu
3zz7KB6Q1nWx/+FFp8RREUQOhp+l7rV1lm6mCZmWcwp+cBB6HC1XG+egqKyYPd2DrCELBK78XDv6
4OkiF/qgASLsgJKKZGn4EnLFL4CwRplmECQN8WabKQIH0F9GxU5vPG9VpZfTaphoX1eoQTz5+m/5
W0Ew8JIMDKD8uT5qbiyHjArxpnTVuPPzBYjPQ3R+7cHZXGPxw5SKlM7Fa17q+S4AzYErrt4YzZpF
YY0fWwNz1Xjid5JozRNC364cXZPssqn8mdjht8/5SPCnHyBBTzhFfgKj2ZPDr8LRj9Fhlx4mZshP
7fJO7wnqf6EAVB8D1zNMatTlvwZg/Q4A99LthLPJoZXNJDX4zn+Cgldpbu31QL9HPGNY7CkOYAJ5
M/55ULbS99KQK6H9rK3L2e+lKSAR6jwYuoRillBN//qLj+ilkVEQ9s8B/rRXxOF9aOZ0beYTHEaF
DSCx1VrSFTpNByB2+MQ9T3p80WuFbkz0L5WqlYy0NGd/pF+oV5mZCZeNJlfZYUixYOqhSxG8bino
pEgFXOM8OGQbM1uZh+jbv/qV5At6HjU663TMR6hQ8e65WJFY54wNYVxQ/9XgWGtxSPebLfP3PKMD
guk6OMF9l+s8OMcoR7CoS9ox5NXaP7wbpX/zbaIEMXjrGRam+L9P2DEGWAc19pN+5XlstXEvKVyj
ehKrMhndC1AnSnk2PPndRVY9fmpZJIA6dEhJhNuNDx9NEu3GYlrjsSoX1sriWMj0IxEq9HJdmfzT
Tv1mgEfZbFPxIE2J9eVeQ1W2FoUlhWInUuTwl51PkniWFP/yzDmsZl6ubBBVFmhvV8b9kcOSa+bk
Ghc+lipBEhbRU5FkLIbloF0YUl5AsntanZp82GFikgoz3FL39yPHEZIcMvyHzFHqayhjThB1lF4K
aL/O/bT6+eZ4s4h8TcHvfCFCZ7NU+dOOjyDfNI7/wFW9dyV6IGU/1n6lCSIaPikjBGGxddAhhVJI
cnq8+te/AivtD2+WJRiU0k7XvuGcCFMMD8PhMPGPhJySDHMOUughy/56ev94zpoV+Poa1aVSlDOc
GsOuB1jc/ZyI5+BxIrugfwZ97JzSjdBk4lLPL52yxuh97p4T0LwIXXPWaa5AIjjDd9X62MXBQWG8
Bp/09+zFmvf7RuwtWro91vJ+jjCFdzAh9q4uJgEN2gU/tiWekqSDXOqPm0EikeGEbC/AlQ30W43S
c5OWW1nDLQsxLOtDqnxxWGm1EaP3R2mOI6DnEfQgf3Ay0X1TYdBEOysfIQ9D38Lod4DcXGrkVXrL
wLcRK3HMoshcDMI2afMxX3SWjkIX8GL9NXlLOnrwifPBn4i/j7b6Qnn0QVyEL+bq7XN3UoM9UjMT
ssjObG8yF7KiKapINVevQ32DEYh3iaHSG+JuAoZeE2RvNNaQvXoUlLZTAVu2A08VFt4bsdcjA1Vq
fLtcGEedf5oo1uGAvRpJ1lpySvkrK5VM2LQ2ULUCAccErHfF/PSlqE2vnCXtxTolRqT2DX5Gdugl
F1lU/UhVTZWLYrQUYz71SD2MaygDjXC9LhSgIwFWF2/DNw/pJzPUASD2FJcKvSgbLQNp2uSG8U+q
e/R29bsmRqC6eaoZ6pcKw91wqeyEK0aa4IoFQ/AuiUh6vLgBdtXNsZlJG9hfu1G4w6hWxHd+Qpsm
UKkOfO19MV7byrRcv6q1GqZh63HJQPbidg7tkWOVE6t8Mr8jpHp9NK6br9eyPFapHzjoLgiN2v4/
rJTYwFr0mwRXnux1u8xg4kvKETNeaQdGdb03hJjeUl+b92WhBD0NFCttS80Xdl5YQ7CDNW5Kqy+a
M05OElQiJwQze8X3hQzUuLXNLA18YK3WTvcx1ZrxLNOR25SpHzQwD7/nTNlfFinYSuA0xblAbO+T
8ABxakZrd5SD8aHgvrTRr0bskvwdKOJasD7fZhykR/RGlP5wlTEDM2kUgA3MHSFK6405kNZW2bUx
VZWbRUfxg9WIMkteTW2PZ1YBQn8HADJ5KCTNTl5146lAgj0Iu0lfSlu2u9lCXPyORJZ/TRgDPBhx
ifqhr3R4ZZMp3+fhJzhkS6EpeFtwqJya0eYoSXYl6wnN410d5OwfvAx4Bxn/hQneu0QB4saw5wre
TVTzU/yVYQ9Vr0eAFAgtizs9uDCE87VBtibzYB9cY0tRQj4vSzAu+7v5JuiwcLeK5fhUU72tmR+i
+nazIT95AiuuB93I34DoLmyLhgRqNzFvXEgb0yGKbzBQ5nMYMJQWZ++bKFNVu/UExr2DYRqAwtvD
UAlUxkIDdGZzyeLYV3GRaGcdWzx8QKQTDDyrt7A7X0zuhmi07WyYnAU83V+nAOfSTUOsOrF6gfrS
CGznD1PC0M24VEMjbAJ7EOp7rrUuKJBXrEY42vwK4q9kSPVd+Fx8dQcfb+ew0kE2WhJB7QfpWJdw
VcKXtAEen4e33v42LJkPaFLa7dIVbQeAbit+3Xlq8+yDQb8a0pQm7vYlAqY441crqL/IUSdy1vk9
p1mvtNby+DhdckbY1PNDvdtjzePTrXAvYMnkELSVYFJtgmOCVlQ4uPq1J8z9E/5TGz0KnHvPAiAR
CNnUeAMM0QGIoiJnA6I/ajoiG5sRrgxESa2WgHqV9EYsM2Ixs/5KWn9nbjZyfkx0e2/Co0rCp2gs
g2kOWNApQQp9yiakF9TtxNpW0V5NfcIUpQF+bvWSFBF6qXPnz22yrjzFipJvVHV+SOHD4UY1JcmB
5q1vEvzAeE6BNS6ICh002qSwU4JtC8ht3qH44QaRVI/oFXJIeZ7t0b1P9w7OiImZ+BNun+kyK2cn
66R7vS7QH0aH3aAqzMA3k85C8SKAgTGIXc++uAZHWFQobpc/CU4s/i7wWAw6gmunB+5T6BPmoiYi
Ds+XnRwcIUNgliQdaauisOL/zOPwZGNjg8e9HOIpyvLxdBSeHklosF9uBrjpcSvETUtReyYCdRpY
2pN1xmFaEfogB7o194GNd5gh8uNHSdln4jLhHClUBAVnuvbSivRZ0RxhWUL0XG7dU0VdKZkfQmtg
D1opAasZNyEHdWcZEJEwglFJLMquUBJjL1t5V0OgGXtMl+zcwNISRVzEa4CUubgwSeE9JtnmEJZY
43YP1jJmZnuSU9jA8x2VkGlMMSM5n7j0jWBuzuwpsx0C7PYnF10WT/QkNbWKuwUXLd7aPNFU4eDg
hm8a7mF55RjQw/x0H2V7ONWMB4dfGQOW23I6HPmV3Nt9KujaNODo3ZeCyplkvWSRpTapIaLqKdjY
Trr0uqy76WBJYKUbwpR/Ahz4aidCvUNBQ/QnEC4CSIQGRIOF9vpwDizLAHt/hr2ZF5yRG4qhGJlZ
ANIEdgHvjCOR1uADMAx4yoW42ILXx4tzYpL8hOgDsR1YPvM6spM6wIRdkPimDcDaUfec3GJc/agW
l1XijpceZM10SbH91k/WFKTa/RckEl/MjrZFXUl55S7RFEFBW3r32nqkSw/fDA/boV+Be/FLwwrY
Fgb+vGnsQk2XejK0qgwjYSzOi5/dJ/BjdK7zLvRbf03wW3Aa0GWRnOwi5RHhqc+/RhS3LnlWfJpe
B4GmHuFl1tu3UijjxJRVZUl8e02qHtYg9BrZ2zSb9wyBEOrWNhRO5Im8mLbVzs9bYPed/f1FAlhb
YcRqnrX7JED4T8dJWep6gwaGKj4uoG9JyPRjQjobYhiP4kknB/inhdU1mUoI3LL7RzeZrNl/E9KG
q3PLxCyD2p+zPdog3/8NsBTLiuOSowK32o3HOWIVe3NQIAMbkU8XFKLv5KbkqO7RR1WXwiuieABn
cfVtLcerb8GMqNBbr+i+4iJaxYqZxz6kyAGzezGtmnnMRPn9MeZRzqjQKJ5/uqRW/cDTLnWWbR1I
dv8HWeeNNo2+EBTzixWarrompk5oSEW6a89GopmzlDsrKEJ3ApUk2mKgPtaCy7nPW58DuaMlUfSq
NhAb7nS81YgaMgMGMWV/jpja53jbjVx6eFIGRw3772ixMDOopqTLPTGoo7zTmXzW3n3WDm91YDnq
2l2brz1inhlDdq+tsOdATXax3gRHt/5x9ZhcRElfov08Yx3HU+7JnJpKtJMuz2iWm7TBzrKPAdKb
163SExVSeT7zsjLSlhx7Fd23Wg2VQnBuXJ7Kl6K2Z4FFKDGxB7bauPBJrJnn/lB5/DFBSyUX7u9V
AWQwRfpjuKWHOrShZ6OBApFnC6i/+Re3qfyNUe1H/UVtKq5fvDSNySU6TCvCdcG35R5JuzCxN8dI
1vszdflf9HhXlXYRb6kYYnoMwb1P4LOv175+XFXV8gjpbMOyFUMK7sL/8KAEbdwB3brPzqqNDjBl
Uwprnz2EgOed2OosN8EgzYdMoss5WcDPZ44hASZdz0R86Kmba8aaZdJzQouQEVZ+AxdOPzveUkx1
ubGmBqQF6al9lHRC8Yq2f3w/ZKSARgy4CJ7qWTrxbxpTnufn+TEutyar8J07AM72VszGB2nqAv+h
5eHFua4gO0NxIaSWEd/eaXudrbUN9VTRc0FAklMGALdEkokDyMARPYLiBeY3jelJJzkuQiI2ECcR
fhXQaNWUc0rX3ipLAZ9xiHcmVZUISXdGPEuEOgYET58hGtfNygowfYzODy5lgO0BHMauEEeHDG5M
M3wHVK7iNgiZCtoX+SBAQf08XriVSYZScFFy2okGjPcE9yv/r993nC2LPfFiuGm+JE9/n/VBRr2n
RHRvxyUthYPQxPet0emuEF3dnJZXj/NAmfWy/NJvt6PK8brlcMCzbfU4kC8MnE/4601tdrzO5vCf
28jUpiggkQv+SvB6Ox0NX35Uwfj1ESnrBEaEwj5Hvkal9v/b2jG9zrKL+Y/TNeVXDdeHr/mpbeFU
Ctmnl1K+rnY0J9hykw+tM6apOBGgwsGrhHEnZ2nHlBjaTCIkoP5U+BevAIrlQT3sN4RNUY+/LO/e
MnpM2cj1xdWdRIjMX7j/lIkSDQXAtC/Ehh5H7u7hIDwqO0HyTDvhQwu4NF8jI9wYwAoeL1QHbxhi
D7+75JIcV+kbgK+l+umOaI4fsdaJYsrhDosxCwZE57i/QsmpGam/qxBrPDS0N3htg6IPbKk5722B
rb16ih+rDyKpfvmlC56wsC0Kumz4ZC7CpDkHHdPHSwkRVEddOsfKx8JKSsOSMlWeRz4gI+U/wny2
b0lbh0VyzfQthj2Rvr3/SyFeEF1GL5YbFfvYtblrAIUz6XM7wm/yVSf9767Opn6ak9ypzfLyo6jX
xo+uKWqbwcOYj4J0r0VY0gK1QgQ0OIKrDBOy44Szr05q8vW/kRaQyYHw6etYeR9gfxHsVEFJmg27
Fo005QnPZYbyxTMa7njF+9cX51wPvywavpvjOYJKcySXqEjtIRiYjK/iVHTL+XjStaP0k+QRd5W0
MTynihFfFKVD7DzvLpj6dygxbjVU8eWyhDJE6PbiNZKiEJ/JHtzhTgewFWHdoNMuMO8YGGfNfYFP
9uh5mri4qPaOzmT1YmAyaL0HiOy7lrKGL/m/+XS6bLNV+6jXYzdnE9OKcDHI8I6v+ILUaoZViTPB
LgNa+UklLaDvdQ6DN0+ImmoQP361fcwEhbGk6E8Lu4nY7GyJ4519sUQcqiS9Fekrxhphn8AL5BeJ
+zYi1mN1v0MQzZt3F+ez+tzSUyZSYeO8fkK9YHxidtWMoZgxF8PCMerDxj5z+sjXTwTEDRcUqeO5
c5znushGztV3zZWU1GBih6teT+CUGUYMPPFgZYb2Q4/Ey73xtzEWlz/8Rt84AY7be74PPoBn9X+o
X/bMFtDm2nt5WRA139bkKFrQOOovhZbFM2/+PcoBtDsT3ypLqwPLY3Ri+hCfHjpaLQW4VhJk0Gs/
Y6MHjnKEcM9VKBJf28ykMihxg6yjhtr9EP+6AqUqu0xlnrA3XcU9ZBSD/tTiI6j+LrNGV/ziH9ii
WHXeRoG5HrdnuUNpuJkyjU7eWHdFY5K82hHdV7YZ4EI0RVNeyP50we6IBrXQNGC7xOnulvM27/3N
SZz+PemhCLEHtdSobHiqYK21sVXQoY/MCulhVQm3rsNnWMC9u75V+gUPqxnOXVgYKhaWzQV/3dTQ
9clm1qiUwgoo1J6Yu2buvQu9qim7LtbkCKpG9eSidUenfVNJJLdoVHgWN7k3ZQjKeWzn8gzn+j7S
/sWD7JCjsOU8D52jc5W1XczAw3kVBIWIwobO3vYRrpJUnuklBk9NPAAVEwDz6/brGbFwcrF7krM9
b4VWV7viAX44sKex2l1ZldBiZuNMPfDydzSqZMZFjzQKYg3Fgv5NmPyf3cND9B/u911WFM2OfjcV
YGuhwryTLjVycmpEzx3w8BY/B5zClJyJN1sKx5kHNk7LoB8qc9qbpCQY+ckYGaMwU8kDPWKQAmwn
Nbw8tranrKMOj6epbu+dOgY8IhPwSTvMpjD5L9l4KQIfBacA46fPb5rpN77G9OsRAR6ZxXfaDQr8
7w3ChifjZuEIt6UZcDKl2sN9KzNXdTmkeu9betRpaO+uRAMsBnaLCLbP0dGSRX+DrXbavEGygOn+
umOzPsmXlNVzab9Db+Kwr/jkyb9QdKhVxGijXrB8oToik3uGRbSIELvuh4JSWSE8I+qEef6Mmhb5
vSuavJQsRhCC0V5ix2sVfFlWTsM9dygyLyRWuv53N3X2RUbEH/tXzgQiWtQBbJkXQmvhu2RwoIxc
ewQyz7ykpjcKzZjSX+CwOWdVfe7RrtWBOabi5fOfga1GL+o3V/fRxybjBpEiU7zeHg4oWxzgnlYm
RVstYcCySGRx+0kLOECXe45QeoejD6l32k+rfFkxGnJQmHYWS+pfzwR8uJLkJTWC1q0Dg8qcsLwC
UuXhJzXnx5BTcVhmjXXgoW1q3jAXI38DMGWLRcjttkLCnVtJqqHPUoC83BGS+8JAOsjH4MhQjT5m
KmkO2qqBBiIOayTyQzV+mU3SLKsJ9UEhPyRPz5yFb7zStIEtBmSQIRVk9m/bMmpZIev30ujAkTgx
O3YUInbUlr+FpkGrNNzWsVUwBj0QH1EIvSqfx9JMcIBVeN247Q/4E5WYXnLnpSlnRlcJCLQ3AGJX
mtIvWfZrZG4hm8HVxLWH1W0rfSm4q2kcinE3dZt3vuRqmgSdDruZyLtnnIUUbBtQZABtITlRqeFO
rYlWlj9KkQPyFrBSkafRtjSa5ekfUUwh6/2NC88SE9nGKyeuejDphBylRciD4Ygz9xLIHUe98+7U
4EF8kxg9mZJg3lFBB0D4riO/4WjTDHWGcFYnbDv79acj43ni3oILNDHxUhM/V1o8ksqUh4F44Egx
LFVnrFRHACwabG+8ngRYuR64QJ5JT9C8q3rDJhQQ5sdrov52w0IxqObfSsGtLbRsN1uRY+miZWmO
x4x+iAtLI33xYBR+24i58EcxeZcmjc6b5J5DU9Ogm4iL0E45vOSrbVL8x5xSiz3+8aHcZtD+dmi3
NNs0w+J0jWU24XlrdcRsCPJMiiSyNPIYisJvrfgcd54RcaqidOnwsBErL+w4lC9rU/7myQ2bXzYd
nJqBG57kT9TTF4otMzO/4NhrTWggd7RRGsgYcfa7bA9WLmIsvPU0SSsd48WybAnnDPdsUHJnh7x+
7K+gtOl1UoJZebalVnHgYB4QuVmOQSocemol4eqxDp0TPONTfc8xWf2X8I/QohDlNF8eXFoEFIAq
hqGPK9Us6Emj5XqzOifubch3yqOkP1sVXaVnFzEEfHk+fF2xsnGblipUlHONuBe/USLY6CF2kdvz
cyPT8QNftGYXQ/XO5kpfYDETHV07c3bzlT+tqM19eelHv45ULMLdNnI41W3WSSLqZoUP/bayF8JK
NFkOJvcKWk5FFrXd358myo1LKqOU89YEFr6ll4v9ZsxiJ0Gxym6XkBquv7SgIAPIDFCdBZqIT0nM
ShGzGqfp3HRaSfq3DiwpvASzwplzGWYIT7lJdXj7USF10W2EpikB+1sgvaxRbUyEYvHQiNdfq92i
/U131tO+UnAC8vBMgaa6qedbXDC8vdO6MvFtZkRETNWqFz2taXPO5/4keejECCNSZAZAKfqubpL2
VmdTSinHa9TkK7O4zX5BXTgsg95SA1Gy/IShcxiJ1ZrAv3x3D/YwppLWIxjnmAkCloS6SdaG5rhk
5hvv+zxa8xM53XCwd13Chvf913ud39qxT3hw37e1xfV6uQIlE16aH/rW+6szuZyTacM8JETWs4A6
rcvGMsHE3tSBg/QBrOeya806YVLkFEzdUGNZccDzBTaDUvR2p/9ssy4ISEey0wIjWCoT4gErd/ia
QsLxNvsRX8LDb7wYNZdV5RFYpph3tqck97R0qEb4Su+rG4WhG43xWkohBdrqayqjajOqdXybwW78
74b6Knv2oF80xaIJBuMTwKMsRyynQM4QZnp3vkhtl4ftbr2M7ZydOTfXBUx27CHlv/H6TF0SFuWJ
I8akhNrQokTC/Eud69J1s1NyIkGrq8M63/fXC6pcVcqtP5hcUU/IE7M/QWc06vuo6TO7t8Ig3T//
r0IUexugfZiocinuu+nkNLC3WKgBeNMB9mOpnMWa6/WmaEPb7gemwKF+tRrR5oJJIl6Cc+doDXNk
nLkox4fBM4bKa3g0lX4tGJQYUpGkmy6uFWl7/Lvq05bmu3lOUZnwfteeVgd94fY0K4FFUR24cwI0
hc8sDuu9gU+NXjlu7aj3c8FMyoeqMpGRgD22+jMbNvFf/sCKcpJQqOdJpBJXa/cE4oV4zqrziIFV
+NJWhOFXlQZ2tCcCM7W+t/Jyqm69UNYCiQuCL2X2V8C9gcTx/Fagh5R8HDx5PTMg5MY8uNzpw7/T
5EFk7iFk4aNlHWFaPQdf0HEMMSLHjlsyL/29hn6LKeNRsCM1HM+YHXBu8oUWuEWQirmaCGnUCUuy
MkmWCXS+deHYyspTB+g1HICCiMGskItlvjbYQlxozIZGJFjoXP1AXOusMFKzrm0uU8UsNBlusB4J
7R+cjQCWR+8OIxcSf4u2xui6pqOu91TebwabSeE2DA5iwT5jxfntunqLuOBAYeIfqomU3CI/Jf+d
vZ2CkwmSTIMD4tbskc64Ba3R7X3dmnapYrXoWieMXZ9Wrr5u281Iuc8kCb6niZlCY2gYl1GlTR8Z
75dQdC/yKOkJ7iK3y7NlHZRV3UMMj67Ko/RM6GtAIXz3eKJ6OMgkCLY1Szx+4vjeJ/+MIxP9pm/w
8csIIWkl92nL5RHVmPCyu3xzfB8MSpmq1tWvVJDqpCX+iJzzaR96V47j35WEmr0xP7mljxwaxkz4
0dhEf3ElwqLQYlF6oVSLP8e4P9mm1bCh40+T28SGWwDqpVtN+1bSmhwNN+c/UvAK+8t2eqhH8BGo
qIDwT/q5ljCpZ+MghWhkteqQl1CKdJ2FOz4MhDG0Q9mSzGt1Nd1uMG2ug2EPdF2PFVMQ22M4WfQK
5rSqTdo47dfzf+BIrBvB1aVeXdA47bMP2sbOhDXkAG9iQF0aT3scxSU+IS0tVc0m2nxuDswAa8cT
62DwLq5Yq2OJu7GIBb0yWnEbmDhIGHfDZjElM7VbpIEcXOctn2EbDis/rUpxZWAO6St0tBziLv8s
vZuorfgXwEM7W+v3l6z0y8ghALGesk6+P02jn2YX/omLeLOeUUHNXmtp1oejYgTkd8N7QLm0pwf8
bzEff9WNX+r7u4eQ1bAQAec3akO+HFoPuwa6lRS2giye5wbHpJP2HegRZ2HA8McVOUm1DOxrFn+d
dePWuep3Lxh4mxYE45gk5kqk2Zd1wnk1k+RgVUqEUWkmqZJhMa8O9NFp7RPeYxRp+QJXhvOKN7R7
nPP6KXKHdyb02CAwXMadjEZs4lMdyNZuoSkwtO9A+6cNebZvJaXGvoH9pZcKYFaclSF41kYeKeio
qhS+crKfqkJO97ucRFLC8TYIV5i+SOtXw5rfDQJJwkrpL+ytLmK/4lMFCM4qMEP/VQZA56Z2HIWq
YmA32sEzEBFEbWHJRMnn6wIFWyzsptJdxdI8PKbnT1rC6okm2k3wSTZzKacpPQcIQRyfvp4maCzy
jBRqaPnM+xiA4Hvge1AbkSngQ38Im0GsuBHO1FaHKntEUAsGv7IsULoyqYfuJ4/G6IhB0f6/3rVb
u1Khi3bQPoCPozja1hxbsZ/MU2lRqRfeO6cpI+5uyDFP+hHAx5otV1k2T3m7ck4ysvctg7mzXWs6
PpAS4CblN7vrASQrQ9H4Kw4mN7wXM+mI4BLidYFr5zusSPywQQaZSFGwP/tXoaHfnbSzbFyIpCxt
B2jGjvhPNSel7HMJPeNKMlocGP8gYOBD+YqBQwCHVO8tF+5cNPcwbqS/PoxmEhIDju+SpGYgbvoJ
WCHscZaak84VSpjK70G761YGC3XcmNvRCp+HtdJoaZlaF3WeqPi2NEd4uiTi6TDJR42qAbnnyvkZ
2p0w0NmyWkJ33eLiWH9rjvCj8y7aNYNmg/YfuH0qnP1S3imPGOb5eyvemZVQ84i4l5gRv4FRPgVU
tgM0+tR9mhc0XDeCEBwKuoD27XKkQD+we0snJ1UX9fftG0y+pxmx5IYU6wjt1vVdm/6LVwoPUpvZ
97eBKV6lJlSlj5ZI9ClEq7ch8ww04KO7jVljAH1OPsHVya6aJ+E5XG0Td5ccuOy0X8P2Zvs1TUjj
JsYasntd0QSuXKMkKQYrzewFJj2XxAF7pI8nGTJDAbeOzq1vWTKhLRDmUsHPk9TB9HEepUMVbi1m
r5mOFqD7ZDxRpu4YD3suJy4J1gA8K24naAxDAIVYxehU0f4sY3egYuDqzehTGQQMwXrYyD2TTcVu
Q9XJyooEZrtrJNp1415poukdboTEfgXGbzpJpNdj5VrCx0ARb5O7u0UkkP+N4ymFGTeGpJHRNrBB
X1S8O+JtqoLo8XtMuWz1Wnn0AlhIM8FCFlncIp8ShwYNxtWJ9sepPbZUlWx+vOdaBSuOysLnwWkL
OrMIunn/632XPo6RChGMR4oWPKHapojSETP2xOYl6mU0TMrbmaoZZser9l6sJFwEKqiBRB6wccgu
Zh6MdSuPk3ijqJa+lKY9Aheau9HL4pFqsTL27Oh//GqsSWDdzGYAZOX3wlnhVrd+8+nQdc2GLoKK
DLiWDC11i+3/JTnUXfwgS1VT2m/rouq2XjBb6icgtRuOMilFVMoi2zspfAeyBoT83QB/xiyBLBPr
D+apltRtxuUfer1rlnMkd2NPMZqAeLLSibCHdjEhpZVBG2w8Lix0fUChJIMuffWGOXaZGkjYkix6
ywN3x2E0gGnNjTSfer5S9/vODLVznL4f8NfSCXtJzpathMtsJZ4xv2PepvUjK5t5weE8pqBUTI3K
ZsBFXDn6lbTcInjmYGiHfaZlnbr3b/JSwFTV77AGQGVAv/ACBLM6+jZjZ1bAvSyIVBLhmLGECDGx
i2wwRfHc1+dBYJ+l7daPfZP4wGCOYHe4BYFGoJM25Mz/frX+K88YadW4uvlZUdpWNWpp2TcRS/t7
XW6QNYczgEHWk+bJxsPs8sn+yYd1NrhBZm8kNWa+ZI1y05gUfKEiFw/fXmDevbQb2dydb/0U7rXJ
yncSG8dNkQ67dK29TM6j0G95zE2sVmRLEKWDFRfrMKuWmrUtyTvjl4TBnEQth0BmPrENg4e4KEdq
d/L3zHEPqm3sQilqYYi1qUI5CQWEYI+ZIGMUIPh5k5kwEwBBMdM3Yc76g83ybeqNGmt+mEV8iv2e
UPgtOVopkizow0+yHEPSKJ0quQj0bcRn+4zXn88iNx3poadaoHmgWRJ4ZouuzK5fFSLG83+4MWX4
+OIyskWswr8FzjQ59AvhxvfTiTLfZr7EuqXyDE6ddBYNFOhrJSC+RHjfH5UZJjhceq4ytYjL3kRX
zOM40b8dyJZmyGbwLIkPhiafUHkNVHcBDLSsEmCLjIHyjeGOiSUsFx5tkDcO5Op/eMLfGJAoAkig
0ZVctt1dGFgcxfhU0EzUpP1ydu7TLeSmJGZbO0HM2Fo+UD23G9dQdJNxU1Sme7cRNnk3igOE6q4m
H9roayWP0h5dBF4Cp5+3nYJX7xWNxglxSCnHrgiu3FfNRdah4urd/Fx8xK3UVTEhXLn4H6NGz2d0
gwEjdmp+TN8QALTlqq0RGdzFUBlBOpqLilX8t3/fo96GGfn0p4nl7w9lP+p5M4ZCOQFXG7FdlVeI
oSvkj9CRV+rtd7mgjviqdfKyleVdLgoGfFhvUOhxkEM+Hay84RRhche+lcXtJif3TENMxrwCC7cj
csk1axuNE6OeiyJBjncbwz/bNUfeD448QQ3wJsKuuoMBoJjNB+8iNNVI81Uii2gw1VyE1JKyptoU
7qy2O69ORY593Bu6l2s3Y3Fkyh/6txlLTFQhCJjJpLiB1soseh9BnQuVXAi6YKemkH2LzsbTrLFJ
Gf1ATab5F9n9/xGZTB7ckimqYabYXDEXCuHbzzUzgLtlsl/GfVd5Kw11HodzwiaWg7PIFP2zUpRj
PDeX6Aa7nKaBLoiRzC5T7s+V7dtUAN6Fmub+JxPCSNR04j1pTewQC0tEnd/MzzeVA/JEIO2NwUhN
k8M56rxxvlDwOBTQAO9at9PMpjjkzMzXELtoKc4gqgDWYfQq2beyH6mC2y4tZKtVCvqH5EsTirw+
oB6h3aUZjz4SFJ4dZsigrreHcrZby1VPy+IaRRO1m4Vkm18ImcUKektZTbKRJejNrXf/QuNpaRi8
45k7iw5k5p1GW8zFHGRcfUmJLHdYNFEV8HftmMvhGSFQx58gsJ3PCuO47KSWyyVq/AXWa8bLaDoV
/MAhhCrBS4WynehJwgy5NdDisW7Xvwy/li5s9WsvOnDjtqYoN4RJwubmvJABrJBp2n9sc5dvZq9X
ZIGC4wGw4tM0SWzwMIwv4+ogy01RHGDl3Om4FNJOLL7aaYX6TL0kmHtFl1yYae9P08c7A8YYfEEH
XeNMrdonzDzWM0/VLnofklBfSuoT+ZbjSEjfdR9aBvahpoK3RwS3g5hqgq24qTF1f19+a/jJ/CU7
BG2taUqZXb70X4HlTe+P86Iy1+wBXCdd0SzNN2dlt7X46hsxJUByGOPbWzakFZ3Qdk+/rr1zyEKV
LZvmMnpj7W2xVvvLw/zxDbbvH8guSnkxVmhZQ1BQ0Y0/8E7yK1fWTlG5S+zr8POZN6DsUvt482Ta
ktl34q7yE71/NJSIxCVIvwHKEg/M5FL0qZ2i2FAedy1kyEdFw2kL9f/0cBULKY3ytEpl0juBjAj4
3QtjsY3BZVNZjucapobO+tAE3Ne4cGKocrRNSvtCJMfBs8LHuFQugCxANhXPrtPjYbkmFo7Z6fu3
0unrB1D/H5YKcXaXtVbeGmilgK3eTo5Abxly3N4iT2u8ITCKMunPi5bGF8UiXTkxM+jQqayE3Tzs
5Dok6E7sGMcDBwxE1tp72GoDQ7QE2oUp8gkZiu62CKh+LHBYsfScMj06OErjbmnrR2/9J8BPw+92
r1MnZK5mAH/PAE62dAnbSW4V8ouF63dMKUQQ3YZTOqgt/B/7M8oSydpCzaI9zrIhGQcdwNJd6QrV
lRCe4cfSTdjKXVHuUr7EV7TPvECxVYSv5m2ZdNWGv/fnQ26OHwo7ruHtd2BE+jlWMc/u2gFygOlr
TFcRLTUxmMskMp1SHuswpp5Yu8md3b20qho/G3V16XTk/EtKYRs/RCDNlv1RxaPHMXrssVu15FJF
Mvs/+13JuElCgreRtf98p12OIrPNAPOBNWOXyd8eQvSIOfl+pgjPslvO2kAk53OYficBJ2YeyY6e
WC5K8mZ6bNrHIOL3UUxyfKJF1VE9W4UFxA46fCSKXansbx+FLxUcsmuSPYyjNTqlCOGDz7MvGGcX
cv5iFQP1CMeI8UtVzEeRFvjzNsiaJWcBdUmWYlokOzB+eCgrC9B3JTiW9ilQw9p9Ph49yvxWp3kZ
p+LWTvwmQzW/moYXqGUeDLf39FOrVo2QbrHiefKSyiYUJuFdVEnpsz15W540eqzE6zoMIl9bed1g
v2Pt9MQcxpWNHC73oDSt2MW3jHCoKXHuIVx7b8l50YvKSdm5WChyZ7W7z2gkALk0gSTqPdgpJA7B
X7QZsrmdteH/cqvHBbf6EXA8lwuGuYjv+S6OAecEYezA+I/FbnUXMY9EO7q3gaPHon6h8S9b7Ld5
hRXrHxMOmlNWNl70DZ6BLr45FeVi4ahBpbrHVX9SR9O7yzuzW+cwHfv3PyJOgJSP1coNPSYZFaLF
5HSkugizqIcZxBWydYEYlC36Y8oPkzx2do/2xs4riUfTmzN4JVyJeLLc2MTX89d8jeu8uKWoV4kF
YI/+FJi88nBq6vDWZ6lcjinD2/igkns+MdHBIRz9As5hsTxRt3KiyvUjH2jYF7h+rOy8LBBkJe7t
iTjU8u7pCwO/1PR9PRwUIOO+dRZwnsRhe8Fm7KHb4CJNi4p++uMyyhj98biE0g1XhK94AWEUlh6l
x6baevEk9/YqifzNQkAvHqOmmWvGsoL0LQk2LktAQHxFmeKZHcuUXAAqJs994MRg38AM33Zh+RmX
Ax84wCKLswj9SK3dPhCUAbdyJCNPpZPQ3X3R8dV1Lk+MUgbXWUr/U9m+z9jXaJu/p6tIXIkRUuMP
knL4rpAtUzc2YRdJKG3bqbgOcwVFDGJVs0qTB3wDz1df/G4jIvdPSKjVx2Fnq4KPtynEpLn1i9lv
ued5xtq3X7kreJoPsCBROUTM8pT1PBPRBA+BSR0tG0kqk05Skf0Z5q9rDrAkzNhkWHT6o64PAqmX
P3WT6arOvQl5KTYqDOJm+Hk+27ODB8Gfmk7YRzkdAHcFFjKn3wuWuLHNsEM4k5WIDDUDBQJwtDzI
9kYMecQaQxRjdOlDifl+xaDPVfKY0tJvvPXdrcbCa1smxjyIFG0hKvnqxLp0Od8Zc0/3iRmx8yEL
8IWFHOCzqlIIsB+vGn9MK2Wc5ByFNKKaxGf0s+M0Y6ul6tTo1FiKHarsJu2o7Tq0CRFVa8jK2Fae
TuYJVn69c/CSOaJpQRtdqmRJyB6ilvK1gbp3sjTgvqiz7SLXKaqeMKrAIDrGK7osP9rKtPOuHvpB
0yPNHxEXgTN/oLw+4JamDvnLFgx9arxwqgZTSjR2lB0Jq7sR+zIFeU+d61Sh8lcfsy5KpyfoouQD
vtWq0YStKkVsFbsWPqLa0hkpuCvy9YK73XHd1E/Uj4zQX0Yk1LH1BYKEfaE2CmRE6R2rxClQnkal
spJzBw9Ww/H7MjVrNCC1PV5u584CUmDX8UjepEKQXMD02SmH4fGCwgSGaosJ4oAXb7WDhtWhsyCW
ftLEtAc1GXRb50Kx8z7URNWlvSYskTJ4iKWeVa16h9NvnRSiYco7s675gyabxJk8EIz0ih9iBeXp
Iy05g74Rc/G4mtUoY7PxqlBEe3yvrzCGWJNdobztC+kIDlzGDWV89egWET0T8+qYhJH4+NSrsrFg
QjPDLp96QCaUMa7mFL3jpNsPz3xHOtTVjFTn4hY8faunKWSJBJsUWeVeaw1U45AxsIDtCQj7SmAu
eF02abebmci/TuamsVyoDQr4i/W4yMKHr7t42IPISLlojLq2eHEfm1nLQlDPtBveCWjITq6EnR1l
HZl49JsXxYN2WlR2FNSWzaH1n7WQWJl8SspqBM5xtcBdZYxxSRFLfDkLcWjcyA3e6bb/6ugUmUIT
mIJriUMOiL/uqWxINA3tXWdlW+RGr6a0U1PcmLa+egCAMQiJTEwo0yPKvd4/eqKiUNrEhKQnItKa
x4g4DqgVHPAoNPBKF62JUydeP+WH8ucO21EscIwdWRfysgQI/amyEONEqBSXuPdTank6cPwMXvzF
ZOsiRS+1UeFVLnX9DjuuSl1famEJ43TMhLvHCBqXp1wYsoHS5nNJjXxsfhjJrVFp7N9l3eaz5Av6
+WMOtKv7KDegABBe1gwO28ZCY8TzusSn2jjza43ZExT3B+VRdCqiouH3aj23LhyiFv1JA015y6Ie
b5SSjgrKFAOsU/MiP2u0mMccAKgAxLQH+O7iOk4Df1GGcJVQyE0053m5tIEmpIlsCta6ApNSE73/
egWar6OGWEz2puyJQHrHp+Vpk387aU/h7Q0+ZianNa+6xbP4bDw8nSsmmsWmxfc/Ap3DpEEX7prJ
xPnAvJbcaly/EmJqTr0YB7SKw6SfMfkUS5KS5Ui+c5rzX3AQm27WU89UOp1Ftc6F1DEyihrIlb0v
O8TUFyfjBC62y81maMaHKQi/QNLLQ6qmZwRQvCv/3dDvJHBwsQi/3BB5OT1274j1SEps/uKTMrso
ETEmkeoTy25KH77TFyBJKREIJz6SqQEtntw+hMHL5P3lnuD/h4j29qTqjhFu2BrE4PrYUUwwpHjb
AqoUJERhxKilmNNAEonHGT/u8i8WP/h1V9nTHm11v9DWXf09yCnFMvycG3+XDdU0DSsQ4ngsexPl
nBYKhYLiuke7IYFip0k47YqNSEMmBrSN5AZYnGximW7ShpyOdMmQK5K3qxe3NgtiJKRpCouIfI3S
8ChokSlw1ffZxVYQMrP62+yrVQ2Q4/6+9wMYKwdvaHUTTe2TF10Y/sLNOmN3E0uTblN6ZAOJB0Tm
ktuNkPaVh1H/Bmug/bSy0df+8nAPZ7+olsNVwrVvnvd5rSltmVILX6/jMeHkyLteEH3QgzqFmb81
jgNDlU28SEKJIjSmNX2TwUlo/YusF82hHgUfmG1lkiFUH+SE8McPP8Z0x4KNqsBQixBhR/vF5/BI
gYz5Bj9izIRgM/7bCulXJEtJ/KsrYgx3g01DWDTiWPtWysAbQLrjRu6JclDsx86WBjgyotPrNTLX
q/95uxIX5Y0TeGMN3NxN1bKqVeOerCg6nBT28kErCXcB5VYANLiZwhTTRdZhrgKB/VoanNyZP4vG
9kS+pPrOeP15RPqebktXhk9+qMY1u3inU0BM0a5flc5o4nMj37EhHEyIUnLXckpgDP4zhv0b+/Re
AznqspICOGd13OFOWdz8jShZHPF/J/uRiHJnmeX3KobcyIlMpb3IYoVV2dYgqLc5mlVJkBkEje5L
lQ5wuy5TGgqfUFS7f9XqAY+wq4cQVGmnX7f4iedXhkfmWiry+MuoJJLrFgIZ/bdpqUbODPAGnV9Z
GuY1v/lp6tivQ7CIccKIGJnrcD0fFqUo4tcQ8B4XfglrqOjr9ZoewEsKi10nBNbZ2yaCQ+wZ/LvX
/8qJ94D3OVbuX+z44YW/zhqZ0DSp1wrGM6WNXDghuM8m6KXE1nP7P/QLQHzcCElTCxDAKLbSlCMR
oM6zHOpJgEYpgzv23EPTDHlRMth3kQtVVEVXXuVwxnoqjYDCAzLquSUhBUB4+vU5jCvNAIhIC7AM
wvrHmZra9tk/PDPINLzKsyZs223h0zf7llPjpIP7OWtTZ3UNPTXKJiFyr/dmF4x391BeAHHVguRW
MrdV/5zdUF1Ki6SFb79BwBqae0vjWWTa7FgP32hr66njEgOq1LsVFr25F6jSZ8pkYuHcgL4UC4Uh
AmpYriQAct0JUlOl1zle4C4Yzac3ZdZ+oEU0YKWs9I+IEKDBtlQTm9wz5xDNLQm9IMLV8RQuj5WY
KwV1FJSak8Nx7EnYXAHSne1WXlLiP/6EMkN8tPvtfopPnnyhRcggvvNbB8I/SAxMcvdKwRZoLs7R
TLmT5opx82vWG2yi6tWFFLNQ6XOei4GngmwcjZwXpw6HpaqDB5pk7CuW+Q9f/MHPTnUIlQ4fc5Tm
WFji6uICFIoWDttAMzQtEEvHlLataFeMnFwH2DZPzi9KL9FGRzHD6ZgPu8r9PmQpKZ5QnQT3EaLz
WSIuwuc41n/ipVpY2PZzACoc5VxEdvPmnWF09aQDSvrtI9E18Nte/UTnplLXxXFydradh6mT7CUx
za1g9g2Oo9J+k2Dwuk9M+I+9IFJVZaNYy3W808xAPoEWLRIgrJXd3UdA6gv65DORJmYJQeUl3R3E
EEEpINnS//7T6ZJ7t0+Elj6VkJ7eLQg3PaxLEUImQqtlzcOYQ8/92lmjAPoz6dvUhYiCikcqBOo4
BbMV5RN60AgiMpJlq19QKE06TPkfG0W400aOiZPH1xoXMM/9OaLIuJHQjmn7BvcQEdMCeQbfbmmS
FpYWYJKyk3mCd8RslgxvjEBpKbkWVcg3dLExpzkzy2QscVg9siKkOSZi2dUPX5HsJ83agvj8A13a
ynVaT/8hqxmVsHiSM1EmPumt0E7snTrwVW6fyRsEN+UB5pw3r8CRjeeoBd6Z94tuAxWAAcq8FHly
mQhujzFauHb+P523ftoaAL2vJw2sZPEZNiWdlOAuC1cRYTdFzBOLWPA8PTewkal7716qfdjS0SKN
wf2d2iHa8wYGDnO9Fsx5HG3KZEgFf3VXRiltT0gcTcdTrAv2e198HJx/QHNWBWAqXsmrknCoHr+f
OJgQXRna4gHL+GjHMX/UTijHCMtDzsGl4kwP3szuQBtjUNHhrQ/9Omb7EUbm/kv5XgiuVqZdrvvm
KKBniv4L3g/sVT7i7HGYs7oX0etMJP/VeeeUdK5URn4JYpccURIfTfGC5q/ja9xvl9tYfXCZ8WNU
mVhW5koWGIu50Q4KHnf9bSzz3KVxSIiaipokl8O6IX45l8Wq3rbrA4KiyfFFS3UQOSfEHDsT/B1e
ZdbQGNTsXJq/c9xvMYng2hdhmAD8zumU0QR8KD0HCxIjeBER8A7TCay2/b6kTWLAYYAULeO6j0Zs
U9fUuTwiey/xvKyuPp5zkTcwlGCFijsn36aa3Kr8ZoMxYfzJj4fv4mikLXHL6m1KFXFQ+/kFQUOJ
RsDBvaO3gVHBF93ItAeg/2e28yoFOyq2eLDZriQoD2QwHlUhb21uOwSMw9Nupgd0a/sk2GdsBkSO
skI5IdXtqo4xV+R9u6Nwt5dFec09nkEe+KK2MG0pHGE5RVEm9Fn6DjLZDuxgRZOpwDU0xaOI7rr5
3cxBi1Yt3+WC7URJvuMml5x711GUwpVQ64Ij9Qy/Rs5NmkNe9CW8ISkrsNqmua4RKL6U7dbCBlkI
yAvDWhMkYf7lituzpb1VDL2ITF/bt+hn1SGku8dXSDvAGkVYunyJxHmoNzAXgVVa2313o8Dna6b8
+e0UcjytqHkjxhHTotN4Mje9WaywVL10jRxrWno6JPpIRnajBHhxVljOJWQkhXKHOSCw1obJKt7R
th1+E6xJCGC8Au2waaTmUg6sjGoyhmaflj7eLcBsdZ9NfRub1nj/wm2D5OStn4i7/FJQzL49FQf3
PJxZQDAC4TmVWRlxEvaODUCTTJJ6QQKZ2drUUZqQxdEHCrQ1Ih1MvGwnGmtyyrFK5LdkgmX9uIvh
qnj8FyF3Fw10rhg9Q8mvmc3/L36GWGRVj6HNT4Q3SDDrsjbfPPpek7fAR8hi/jaQDIGJGcbPsSJW
RglUOGfZvmnueaJsqXgAujN/G8Q6t8h13/VC7CHmzETiZ31EQtnFrtKy6hV+FpfWQJvvtObrX1yk
/25Yx+4cRC+hCcwTbh4ekJrIEsWExfuzIjxD9P3BbU11mOKa26uONP0Bnoiq0XQN+CljD7DXNwEQ
xzggoUOpEsGbuMHGoOK6SvKEz5PIB8zFdTTJttPf4dVNnptCL7S4bC2K4KdTLNBrprE6G5384wwA
6FvQoMJ7jn+wpAq8lUTNWCFgjTNIivuz7MGBVqc6oEnKZMbRCXIvIbXiBzwRU+XMQjuBXTrELesd
UoLKSRVKzDhsXjd1hwymYhaBG9iHgf8Z3gXY4hzo+yN4PNplpJ7DDubULCi4LWAZArPsOvo1bT35
LBamTXQHTpsujI3erW7+aZ2QSzifVaCDeiTNgERZSp3RRqdHAgQKiATo3rNopoz5KE3VPotV38DG
UEZEcINwJsI20dqecW5iIR7mKlbHFsbv4oICslbp13UbRjWO3uVEtUWZvwfOvhYtupQnALCl9go7
up4wL1BVQyeu3h0GAqjng59DpPf7xMBcrjtLcCjbzzGf+v17Ety1UQDADt1LwMVUH707hSPt/8eL
oQExH4f7KzX+DM1+Ch2vUSVN6xjz0MJIXcZ4wjKbFWekjfZ09eESCD86NV1eH8ZDHBw4om7sgpiB
ZllaRTgJhiXo90hHCASpi1Fz8PHvHM1t4amIUHS4RLg+t45mVOx6FtDYgHP0894rUhKV/4iKc4Qy
nryIgGuWlkIsbucHOg0hFdLn0m3xwhZGTr4XYqj4Id8C5MQbqBzl6i96YZsgXZK+dvhcQXg4QBf+
IZu27lPXUgLuSAgKhTyLRcJAgVl49KqpTFopBCd91aHdsqznlh9EDkS4qeH9GBKiKUNKSjSMv5cR
qRIxjWA7JqLmt6JwKjfmrqgNXBiwM/UCD35e//93vtGDmMM6GHHyzpAkSyDhapEdjkxcI7DOHUWP
Ex0pt7fAEDNmkc2W2UqQ3lITBIgYA4UjgjaRMP8BY3YrzGsvH5RleNWz9ZQDBZ3Xd6QrlAiED2oe
x8D74ikwLV1Q81TJpndNpzVZLgmfzIGVrh1EVe5HDW1es977Sne0u5dYufZh2+/kHOJSmIh0hcRy
nFT+tbpNEqObMjX+JNHovMhHyBPgfvzAUHbZDOATkKQwdJHuhSaG9DyLDJ/ShOGyD0QK0lHz6Ykw
mLgSgvILKSIPv/crnG4Mhp+HClSl6kgnQe7Er1su+CT5hLd+XJSqicCk6aw+Bq0vEaUGk/GmRpsB
kImNmavBa8R0P8xfuWo1x0C1jg/SIZ54mZO6wM8OmKWecvL1U3vea1VEH8fBuCjfDsYjZMeGRUBE
C0Y/+hogV2aVuUDfITvWQ6i2fdhvjQIgz9sgfOl68eZLK8jHb0sjSqHplw+7o5dKpaOvHICaed8G
a2n2ZFj7aCgwsveAXbhna1GWVWJmMCT+hYcZAtYT5BnyHDkaCcN+iFHfgr8lrontriC6VTsnSbyk
otfBt5lgBFnq5qg2Jocucpm7AcbKjWJgC+aWvN2HAj1DDB7sk+drryaQrcXuTWntx5wv5mipt6aW
4eNs28y58B3ctS6OyEhsFotIj/enF9Ep7bClE3dx+xsRE0Kd4jS1S6HgwL7PFP5x657hEvU2yLqs
XM89sdEz5KmwgJQ9XVq4IfVl8+gIXw/4CCWT65C/26VWB079cygS626I2iPyGL30Ry5G8FtWtZdo
bS7Wf5bH2W7OW+UBh+80ifIaRpm0d29I2J21fiUCk0BpxJ0ZA6VedIrCscZlCsbFOon3TsTU0nda
9XrKVkQKR2AwjOyuQHfXn+FohiR20UF7PYqqDuGJDKAMdgnzi/XiM1RaIKOnykbl68m5kcVUEE0/
BNHVSp2EL7ouZz9kBtHphbLtSB2wxrps3qNHkaXNYeLJOak02VjxOI0tE27pAOAnrCK8n8qMJs6J
bCASHV8JqIrtSRLAr7NKjNt7YhXnBZD2C442GiEcmAZd34+hG9zofyETVBcXROcmWPBcxYqPNe97
81oW799xaYDts2UgXzua7KsxrfKr0u9HqKpRTnbwa4OLIkicJLHmSqZRbNqYqeYtCfipCURrvnpT
w5qQQgrC5U7/BxXPp4hux1qixO8siKnmCbFllhIMBtrm2e/485VHF95F1ga3z0xPmDeP6jbbIQZk
JdMZYMjhfzDbWfcMvhJXiaSRCRBRuiv6ZJEhtBpaxU7kHpSd+9APe8Op5mvvU6JfwnZP0GRAWHc6
hgu4qElJ66wLPiQ9YKNPVw9ZY5kj7+jV+2NW4ryhIiOyoakforuoOEwYGVXD+FTJ8C0X1fJ88BQq
+ZDguGLnTNg/r3ROZwCvYByPZJCyx7yNoalF+1g1tkjKKnU8xxQYnfrXASjSVj8LWpk8pWnsXEyN
pOHpSwuL2oBwUqy3bqLm5XdBnte1MFPTo52pE4bBi4q56ewMjvZ00ADgk4RDSD2TjgqX55NDV9rC
xbWae57vD/Tf82qwZZHEd4JWn1dKjzp9mz27Q6ebEdUtShaOmXYXrmCdzfy9+xm9q8uqfhl74Hid
DgGU+haoKJr9WYfusEG06GY2981VsOUxnK9e3/pdSASz8d+Bwj4txLtZL+TSha2bq4h3/rZDjNYy
WTA5J2GiqTcVzXvbrcFVIaghNWj59OpsY93bP6B2DDsRanSJ9TJxA/HdGTruzMJECshImf1hBszz
b9IrECweBkNlBcTAKBSjyImzOBroWhg6YwuqGERxngifL7Ezk9TeDpaApSABsaUsCIar0HvgqZxU
fsExTQbrD4jrCflkY9liCfgqu/v7Gggd66f8JbSDqXqkV9MchsETYgIqQDSKlfeWw+zmoIC+oCQK
6ODVxwAoHf6EilGXEC0eNK0goUlEf6KXxDWw3G/bAn4aSzxMYr0BKN3be/WfL0Ajsn/EGxrRJ+SP
78dHWyW0Mtix1rTtXjEI1FY7u3+Yaxsnuh4bzWAPaBGR8low2GDvT8XXaAf3hAfmlAZ1iWZJS8KV
V1OaAc59cDqwniOtIPiBWSGtUXQLAODq5/CvQ4u0AJOQeKx6JlxrP5FwgararnWPW3f6lQlWrdGj
S2qFLBQlyfcBKRea5DDQOTRX7kaEn79hLwazcg0kU3TzAloNSLZRHsQ8o0JDa42qiUn1Si3JTw9F
xPs5mP8jQZN/bbEjvWe1jqCyOBvv7wR/UnE4ib0jRNJCyg/Q69oVOnnu4m/DpikkIK0MowefryPJ
DTkPjflSSKnPplZpN0SoU0a1vnM8j7+evTSLHcQsPR0z0h3igKyoTgH1hsqZ5zMQkAYfkV5q6b8X
4H77wLtnBDZ4Uv7eLhNPw/uyo9TCSzpR3+7SmnqHh6SilnsMyBUK7vvGhU5ql3sS4kgGjBEHaAhU
xJ1g14Xr0iCdC+ud7y48Y7wCvp37vXEqc+Jq80bhSSkDLc3NwZ88n+wi/FtDYyuq55JF+2yedpz2
2CV7EMvCzDN8LuWTO9Or9L0M1oOokNOcyhBsq254wdNIxL0x2NxuD4xfdGJjxqerlu4td+xPFSut
9BqbpdGCjFxDRr6FEK5H/LpDNKKZVutKgr3NtMc0G59AxTjAFFeLRfevK9RJalVLtuAGz+2RKY9t
J0npRSU6dD2p+fYLsZ1jy7FNVzXPtw0JITBA+q+GCyfWtidR9zCAIQHgx+QfvWVHZra0A6snY9IL
dyYnOrQtTZvL7WnCNY4WwJt+OecBnKhSFsmzktdYda4wndsz1F2InrvldQ5OEH777uB7eZ+H6uib
bALrluKQ1QClHnaYJ/3KaPoP2YCJPItDsWp8IOYDh1nKJ7ShZAXVVRLy+kKSzd5VIVNkBUJmveIV
GUYaHHSabVTAm4QFcrAFIWQqfLEV4/7Uv3wZyS8w+Ub98c1UdMzs3++/FpIGn70wNtAo0sqd7QJg
CsyOwMZUbDERih9BZZdA46J8gyfVHGAfPm5sjrZkGsSzsDXD2N/n/7UP1vZUOGGrn1jeUSQ6nyqs
uIN6dzsr/WpsHyCptAWNGQzcefNbA4wSexw9WSn0TbMExRunHopbfe8UpDlyhrvwdjYV1ZL/A5zL
/+Df0RWIAn6wSOzbmFETUbD/Z2Ywy2CaUWBpjnIKpHX2EwTCbF3akCTsB+9kKPfjP7rKuxluThrm
4gszWBp6aKDcmrJukjsdUL55RykDsbiKVl1eXI/BqKNK7op+0UipArNVC/MWpHl+k+IeGChayZTz
FuuLEg0wpY8TEi48DEKwmcDB3SHAnmS9PnuEz7nBXwv0FlwnYA8aOStLOtJjeDL2gM9Ob1OZUSxy
MieMTvxDFpQelEkMKkjA90c2fzvwZ4XjsMH67IPqO5zMwl62uJNgDIdB16Vo1Dx5XvZcBzLCu6sG
scBjk1L7Z6UcaFGLpPhLp3fW2Q/lsNenNi1BlOuCXnyiDdUZSyEiOq+dX1FA4bSN4CzkTUkOOo1b
gyZL9eh6u2jsKmYL0QKh5BxtOSDsp1fAVfmg1M6cwxpV2efJafc2gHpVjaF+SguS1FfNuv/vodvm
/zMu3zs6JHWu3E9D4iEtfh4t4ewCfQbgGZ8N9EB2yXtfDDEvEPszhrTih5wxPS3se4IepPR7Xh6c
vRUEvY5e++qobJdZSuji5qFMVV+on1qgfOAx//Bhb8TUyAcnxOm7+vvCSscH57Vm1NZ6CX0hJnFR
wcm4smdWZwZ4/F4bhjBellgDg0NCFdX/K5qvCeAyZP3QwJxBcZuPmiwXEOOTj9vAPbsOhP/EFa1r
txoNnh8blevtXh7aNRZ2ZF56cuAywascvaGZcTlemLamjfzELmG/+eHrgjyY7277fEcuObywbyio
1LbtDF7QRpAeJuEfuHN0zaWFJY5LuhI9WhmmF3YJTDXcVfh9/ZOkeUDFj7UWhQrzMdT3nUr6rOKg
FsmgS/4ZiSinklWPLSVrMW6sj5Qvur2FLbBSzTN0PFAZUrGgV3P0ipZyoIbOiBGD+TXUlcbCmuG9
x1S5JtOaXOB7uHMWvQ8q4DBQqnDwp6ZwP6Z/2CyKkzaZdO5doEskgCxF34gNVJtAO1ZMknk8xVDo
jrUz5dVDV8aaLqjBkMciKEzqypj7ND9U60x6IyW2D777qHZZtg3983FN0KYxxTy9K5xwBWKM3+dY
f99Fd53vLgLXcYyFjlbVpQFJQYZ0oJY7FNZn1FcQUXRV63pmd3/tWUHLb5eWBXIbiQBtHttfDLs4
749f9YmCZWXRUwiBm8aV0vquMIFoxsC3Ap5vDmgXF+SVMJrrIF5x8oCKYc8xfvPBRVM5lzdpnSPZ
BYtfRkcbs9cPwzTsyQPd2Ps9EEENL5lQJRwH5ookdzEN1tG0buoeGHGYGjzxJJ1RdQWuowOul/v1
IetDP4op7IczrSjQDIkQ34I7EOovyChnU8UQ9oaAjnHoqlQ5I/7XVuxAqop2daQHKkuEvlBwuibI
fmqyWjQHWFd6knBQ+FVEmQY+K/5NCRlHEgjYth2d/Sh51GPUu76Kb6cmFXDNG/NpV39KbYBUZqtZ
RrhEFYGgUeV/1nv2nuJYEq030Z7WNWU9j8j5/4/n1qoSZpMh5ir6mU0Ru+g2T7KR8LZUk3RQPUPf
ZKMsc6phNjIZruSBj+jWMkC0SvLk1G8CUV/w26KjM9hPoRw/SEAWGe7b8Y+CI+gR2iCtu0L4H+V5
x06sOADMuPear39sIRr1LfT9ce6A5SLGThHsvT9wNppOA4KTYttpxHFN7KLvgGaul4K2bteMLd9F
5BHI8i4Q4nRiCeliCrAl9FZILUfot2gWwdcCs9HQNIKzjhuam8bjv5SLQrJ0PkcVtrgRYXf0vpUU
wJzMuHXh8eum4Todovikb5s4Df+3xf0s4XhuYQDssusYeD6UCZc2B+9N6zi6kibeMJW391HufU6R
QFRWIvpXU+5pIwMkuwnhHt7D0HXVVMTGQIo3rp6xGa9OxHP0nGGdQWVJIygu5hCRCK9eFV4V86gG
K+nhrncLaWFOxGmm4Pc29AERZN1DS6mRtrnF6BerOTD7vfaDLWR9Xm+yxHPKoWL4Wr2D7KVLYS4D
Tv5J87eI0H2qM5kgxd+892WZE4MI242vP+jko1/EOLp+jo0yjxP9hsiaUOPE4zx2A0/USXNChMNS
Houwo0eJH3r+dBLzlYq9R1x7Em7WZ82iodOu7/bFEBFVDTiWvLdqDfytFPVCm6XzjXx6zltWmD2f
0aTONxaNgGFSCbM0+zwBkztOtqzYkdLMlNmcI6yDh5leziVSNefsDhdbN7g5dnXd4AR4ZvxjX4OW
coHwrngIq/QsRnrkK0q2Y4wAkuYj33Oe7OVCNTHFFeeTXYGOVImQEZKjRSHPBH+nLUipiTMDQX6X
HNqvUKUY4esPy2YcdkzEFLBYfQOxFHpGsd6NU+ynJW3efck6eHdfTLnXAOmDIrzScOs0/Jny8cWd
3vRQ8rNYrRD0ySCdXAHeU+DE9Azxp/nszsMDgZjhWQUWEXAjLc6sAVphhwDLy3Qes+/fJ1FnHeIU
OlnU78/LPOa98YPMnaIK4YzdmW7t4M1F/0MwwiicFRRukTMcZEl0zDHoHeYdfa82KTpsBOjqYOO9
L+k/GJ7Xhd0NZFEGDpfHUM1FBclJ7lPgbyckIwXT8coPTCnwMIPpHkwBNe+8rfqsjj1hzrH9Rb+w
EfLbohcq//hvL+uR6pQNi1exv56gMv289Yr0d1f8lpD/Id+eyFYYtS1q2otH8D/9jOqRCOpN+yUi
g1OeVyWk3E4Gn8C7keIPtwG4ENNvGTqEudkmIaQ3SYDdkf73XIQwHQnskcHSTuCRaQHYA168oEED
mNxK3UMLk1I14yt8FHxN2MKmtrjtLtF/hnT2ez9IDq5vUnD7+PaoH+MZHTCijVtt02qo/NhRum+V
sxCZ1Qb4/ZscPHcDlQV70AVT6DCDR7yLBTTm7WLQIiM9VRRtdzSAhIaD69m7wHRbk99Yfo487OyE
0yZPna1m1xV+jE0Smw//ZAxgzrKafq61igkIn8a1leiH7TQrVfj/v8l5Ly+ZMY4yCHidGx7WyPLN
ZbFb5Vtwly2WzMjOR7SbyOc7d20Qh59QzkxSc7EoTIZ8QeIL0wKiJYTkZI6b7jVpqlSnltD5k5qL
bKC5J8RFIAgd6aF+zAa3ycHrjv4TK0eg97+TCgn6Xc6YFj33MybqoKEa6G0VaBg5QBH6Fx5TVMed
UC1j7E61dgmvKRbRHNKZUqVpVS/viBFfeteDk/7rfyDTw3shKE2jgi6OQ2QPeHvnw/800s+JZv0q
YwW1ukYnQoL4KTjl2LDAwNLc69flXQO5Iq0uv8/pZCHBEvPz5qRjF6IzB3+64ZaucxoRySJDZLeM
AAxB9LDRTpoWsZCewybjRKtLv23ujJTJHIREAsfk3miJRwl4vikn5C6cNoax67sNYl5BYGfV2zK0
EWy/NtF5XpYUngAhfIqJwBO8ZSt4N/sNiISubHbwvijydKmS/pEk8EPEnM6UG41gMI4Az+GqArol
KSgr1VRzHD1hcDSf0/ZMDWmmCuYQRYlewqWdC2wdPEpAnty/BrzZIqUygV7Fa7+s6dBCifi8+B4o
prk7NB5pJiy49nqJvLOavNbrrOFxNmepg0EzdCNlNtvqNIozq7CQoxgfqQ0rEwI5Q0QwOuQEDYIV
ZBzW5FnXSUE5514KVp0Fjig2xlzjxpU2V0hvdAeUjAvE2F+T6L4vOs7VKjM5uNXeVwFEeyea7u1X
uMncykJGDY92ZCWUzAQtwrrDgCSV9ZkhYJrNQ9bNp4UpiBf+Ejnn0LrISDN+vhvOeHwkR7pooUZB
olmIG16/Xzl2yE4zCwDcWc2g2jXpp5RcWhPLjXa+7doDrS+GIctnkASMOj/xIOtL0d+xtDxOKcOK
vTqztcYrrkC5VcGMpWnBfvRJWP2QsBcS3oDSBISwkyagfa44hrTEFNXVT/5tuPlYsTDye4oiITA1
5OBrcwsIM5LdL1rutjxqCFHF1/cLCKtlZ8pq03P5VrX/MMT+yvRT84jbUXI7zrP9DjEgdxanwqrA
Uz879KW+xkkFzIzhf8TgjDRUfjbJJtip+cdfLzpIscaw91TxjY3WpFFqWhd5faV3HRCnGIDJks2N
QuDdjgpNQkP6/htW9ByRXN2j6u9ygKhZOLeTvZAav4MxSsAgSSZgK0n1GQ7nKd2GXDaPLXEt92Qu
2ix0qDyjlrrhdznF/NAc5+cmpCPbSFVEP5aUfNUguEJNv832guV5WqMq8jFwkzoa/8Ge1Zkr2Zv7
Hmw4phZx8LS/R1L/dVMmsX/egzy9r2cu8OEQ5fBwQjsP1y5JZgscofW1JSBNK7XBl1GInkY4xCGA
bJNA03RWrNIAQujmKyHi9qVKHKJJ0Bu3IEgLYyv7k9UfEbnJRoZj4JbGwAnP+nO0xlS4zIuc6Civ
JoDnhqnf5hLvcUBAVxD8JdUqKmY3Dtz5JdpEXCuBQpy3W+vI01XhKYT3gGAKrJf+X9SPIMrGh5F4
4iNyrqt9iSwAINYgMZwWy8oQ2+x/skQcGxas4FTH6lD6BGmDzaxO8YJ5NbrK7h48FJslmCXHb45H
h4BPoalEJySdqFF+xZfG2l25161zOoxn8TZJmB8Hi+Bvvn9A+4xefYaexs7COHNd+ENfR9krJYWD
1JHGEvgGw14wqjndWlBplgitwKJMxRbj/VcqW2jDYl/y6eDzpPuH5qm9XLhmN7cdts8w/f6dr8VG
+MAQJuQyPPAGcnlA7CQHxyx/AcJ2RP2kfBtUWTXYX31/cfb80PK69swmOv7s9MP6yF/o+5jn1xY7
hJ0SpHlSmV8Cq/clFqj0WS6eiNl4YWUyEzme9w2R+jDRQa9dN9dmwg8trpbzn5jQiUsGP+cFNDsV
R4SjdkzeZhEKIOqw1F4QuQWDOM1mIvL4PZZB3PMPWqw9Tw+NxqRwSTUNmEIE4JqSSUzTufJLkTZW
MEVLxhSrrjH9jECcyaG8uEnjsocTnM8/+VjIUhi0FcGSjhgJM9t6ruYqNvmd6BsKa6vJMNIic2XY
AN220T7QuFiLfkXq8D18pPUTTvQ3y+rsvlD7aarE4z8BH5OI0j+DLr8W44rTYVcr2/cgnFnnSihW
gcWbkJIeYWizLv/7NbM130K1jv8G0WZUdZvsh7vxin+SL4pTvIlZz0zRz+ccYSbSlG8d0JvqflAu
nhNWmKYLgnf7N6vBDKEBww8toYc42/pij3cBqfoS47JYFoYNGP0PIN4YqFf7PlM8UORDbnmP9DHu
jHdVc81x9H1oXQuc7Q1blftdQ0kIp2X/g022kGTM2jaVDLgeyfVWjtYH92iWvntreqlvmhrNh519
LxgbwD5otqCOHfCd9Bzd3dNmj1n2S5x/DkH/roNocSEtYjyO6Yt8VDylDE1rghhRVkJNqOl7/CSC
vYik2lIOCSj/u1y8merMfQHMbgV3gSg7PdhBsr+ZqzTAZMBxZG914LjMRdOWUJtiuLbG2PrAvP9o
gtlCEBbkYgYtlLbZv/0lwMnTISbOdJp3kmNM6pWZihjaWgcYqoTDTqkt0IeFF+3JbbvPkZLRAua/
qTUHFMv0EKxUmcj8uXw2YRXRrHpchbUNPsIpT6hBxbUrhcfpil18Bm52LEiROJNpWC5cWeQ5FDUx
XXDtOvajaQYLKSjcZw3Zpkpz7FNrng+6CxTrzNLUQ/KuoDJafN5wKB6jb0oTBNMU5TkMEYjf/BK+
2jDoiuLl2jOCrMHjk4j16ww6dkIsMQW4yD5PAA3RRMm13sX3Il2oAdkEOrCrZn+M1aETDC5sAHTC
30h+sNBS2OamLr1Oksb5p+fShPtiW0soGs2t7pHuwet66XXheZAOkDsRwOlhXooUpKHzZLOwo6YX
SRcZ0RFZmOM22hJvZaLJ27uIfVAwH9bEYF43uJ/iFzZ5yu+TIhPOP+HPAY7mKD77LBncxD7xlvd9
4x9T2zs7LaSfnJgMgS/Yb+3S0ugV7zt3RCbF2D820Y3oIXV8kRNUF2uYDFzq72R7783m2dP8sbTV
x5hXJdxeiedI49qLH0E+aTM4f/r4Gk+l+Bl5AgRxxmjeFNfyu4DTo5tNvNItHu3zOGSWPwqrlYO+
GrJSoulOobFjYbtup2Oz82hkXgPDVwWAEiMELO+ZbxJBImSHrKCXAEVOGt2MJKpVuN5zn3phNs11
OMDny8KtcNKO00rpI5Z7/B3qrz/Q0j3Tt1Hlz6bj1o8HaH6p1QjVeihsPl5HRjnFxZKH1RwJvFXZ
Cug2Ww6V3owhWv4DGuYGTajoThrqSQKQiuAqlm5/NByyMkZANewLPjltG1mGIXgHjL9wDtKuYiA3
u8q4lzP65s4a3sEB/Mq9KUL3LX5MO8ac6SnyDj0a2AVtNIPYtSGJtwuLZJu3gr4MssNYWhx+mR7J
nW1EPnBnsdhm6LhdGDE1AtB80r1mbyI9RZV29C/4xOSCYe6O72bDC7ruGsqOcMivabVDzFbf/8ZA
aQFlEYOctu+7Y74sIW/LKdBPuBAf8kkcuvnRUZTIhl3UmV1toaMDq7rRsMDnrEa+VJtW7o+/q3tm
32h9Wyf72cCX2KDz64rEB+qu/zFchQqbhKmuvbFd5wxKwxHSvk1JntOv3CMi9BpwNuVIAQ9aO1bf
+HhKXDkTjy0ZdnFISnLjnZfYE9ezEE1GWx+tFfvBywpaQM843a8Khyg9rPgYlNGhliq3v/KBw1TE
T/0gY4P34MoKJckxVU29lrBe5KbVLw/R9Vv6QrenTIBy473A27lbG414tf42NQPB/nFbt4kReeDt
8tmctPQJFxdncw3rbMMgKoon0jFmZMOq/4fQZ/j2b3kmXylBcnIG+EQcsyAyPTBFjwTwp4cKWCN+
qIEr5B/ofVdkYHvuTDrIK8AcbgFFDE5CQEd/LopnYpA3/bQTITEE9xi6p40xhCfMWfrqw+HoFIcY
yqlkgGTCbVWiKkqEJMhgAWIltY6cmO88DumtrH/elzKaxz9z1SJhBQ3Z3Hn+gftdJTAJ+7iWVa5O
q4WznBQg1UsF7W+xraz6Ovjtotj7UR5hlGtIRl/U+wTdG3B8TjlL2WN1YUxfku+UZVPjZTuH3OOy
O5O6+aAfnCX5B2yj07Szcr1WVTt+uPhL5XIyrgowZKIxB1afHRi/cb+vThqdy6D3bcPP/HQIrO/S
fMdISZ0F6Y+9xIXS6iTSXQPoy1wGHPEzp5eyaBUERe5Dgvrpq2fm/fPdxIW8BtE7Lt3f4cBMUsww
4hSzZZfhI6rmc/uGCDRTtwLalJDII/2pvZJcG22XCyDc7NwD215s1KPwy5twLXP9/q3Cv/a0ABoh
8mqjpt5Te8Or3HfA1MUpXsr1Z+R7K6eNA+Oe6hUaYEMAExsCrjMDRutBppVQ6214llj2ApqCVbT5
emo2bDdPF+hUufrZVMTtDHkvqIKLRFyuA+e8HJbSf2NUPW/Zu3tyMJl24KPD2u04j0PFWlKeGMoX
npbv0RVUF4sgZOdeVYDcsFFKcbKoMop6TGOR1h+suYlaJLkoaG/iki5ITTNT+AvHLvVLytMvyUXP
6Fwx6NUeGta+cRUnLh+zLfZIw3/QBUo06DSJjMbEjS/fLAcgM7pXf0NChiHIPZuPc3913Qsnab/C
MSHo/+8M2e2Ydh239g5nqyR1EEnAg+9ubQNIenIvH+aZwc2CJFleGLilA+U9bJTHd3rZ43CVh7id
7DQ2nNROiLwn0aL36MN6tkSJgMNCuXK1HyWi7jjby95lEIVd3P6+v7Qj7ueycomzQ89v2LIad/c7
xN8I2npnkJW1G8o3/pEHDRuBnSeCBjlMKPsO0Li+bkcvYXPOouE2Up6u1YARojEhLJo7yrM3LfFT
frrTyapoq6FKWqjLlHQdRXPHQf//QVGtp7ljIe4IC9idvsCIMP4cDFpUKBcbUozOeVBq2dSdmNV7
0IB4zz9Q7myRrW4eosiEubCP24gGZSG/2y664BWwver5+9/8yBl5rOtcV9ArplBooi2g9Gz+XNHB
jK9xm/FcEJrU2MvpkFRzAT2+IFRf5HygjCWD0+j0KZCXD/PFG4JDxQpaZeBmQe2tCE0YSrmboL2U
A/zLSxLEL/rkGdTT93Cqicc59BAitd+JEiqFSdI3YINfAuF1+R/WwErOHK9VxvWHdsalncM4CgbB
ZA6hV7VWDYeSDgMNPmKa8nUsLQyYTsgsggxLDf6cG3cyb18g/2Y+N7mvUF6T9/mpgM5SVsiV/X95
9ISE/gmtLZvq6qdfsKfUt0MTGxNlroujuYHpsH1SxLIck9ifkg/wXSaDvTiP2Os15h5vkStanFSZ
EIb0JBr0BP1t8cHaseEaG7ppwv3rOK8gxfO7dMsXze+QbQTiUx9oiQ4QgmScem+8Mo5ON3ppvfXz
8RM3+HU8+yNjGVx+dJq2kijsh6i7aW8/5O7RkBhaZcBy60aUV/50iCoh0qpgDQJxvQ7i2UAheXZg
aH+ZtR0OepWG54eucPmr6j39tKJ7UcZEtolT3oIQ49L5YKEoZVW26xv1geVHM5FVdnaRP655c3Em
gD0j78SA1OxmRNO+daxRZvgCoFdwvFtMJj3n32tU7iIbXUaZXi8ewMEBYbClgLI27TWgFh/diAnK
1fxgdeBq/dFIlTrB0ppFg62igLg+DLXl/yaI1/T5q5qQN/uwXiE+9mvlkjtFLOPAxG/WwfUDCJbN
IkafLH3wvbFDazdYnzVUiNB83zV2K3FFu4tpKn3Mbctw4npUK/w1TNT5JfthzNFM28yIp8IZQQS2
MOcrqt9YQxpzSplvDHufLHJOj68uiuGjLBJ0QBAsc4NVd9SS1NkUMhv5EZheC3vNxTS75AmPc7MU
oUGByCd+W1wJa4hEUQPwNh3xfGlIecoexmUnx+uQXH5WAf2KDeIO+9112gip4TqCG6dtlj6bf4eq
4IaZ9u8USNJOYKHvbzXyI+z+VMcArOwQ5y/Mx0JgTpCnkU+mvtPi9KvVlg1XAxhkIuO6bIEuBRop
JvaLqJbeZ5CMRv7lCsqpk70GslKvsy+08kHRxGF2WDJrQBHkFNEi7oQoBHgGKq0Hh6VN2BuS184D
l4XNsREO41qmAkq3AwZENcgS7rY+GfHjnJjPnIs6D0rfvV+syq8ASdVBneUed+zPUUJBiYM75eJM
iEJ6KxJYKXW0zOGWKVlFU+sm4Qvqydn+rfFOUjwEQ5vwuxZHoH1I8KUeiScpLe+SzM8Gb18hS1Y9
RvuBTRlqYSdjk4SsubSZK7rMp1ozm+eSjS2xW+gVGPN8z6ccLnGW9MfYdPsuTkaOIUL3gUrai3tc
mf1EoH+jtZeseXSStgztzqkKkGGl3d9Kq1dO6RPgYg3bZbxoFuTw+B+Xfu2rGeRdHaEjJKgmMyy5
3KbDbbOznP2amh/PW1Jcwsfpk+Dei+awygOXzs0Uj4WshYZS5ATzQyooV6nxf6a7aBfOEAPlbf11
eFYKke0FHA76Zz/EydaziPP4nUXZelK3Tky+6d4j/opZ/2rvf2iqHokqS+1pVh4EdRifuLAAEJJ2
vJ8Vox9St/vaYyywRzw3hjptLISv//x/yGN2/8m7496wTkZW4cVpcSxubI+DX8yEqURmFGJ3+yTE
T8TR+TiDW5iL0/XB3d/ZxR+Oiez8w0d0oQTU3qi2k3dwFBgK3RPoAbwZABqMKo8vR5zQN6FsfsP+
iBoHq8b4KVIvJtIugDDaJx1V1WEz7eOIkkKyGvwlsbL0rdd+Z4QMTQ2lQ2KuUtue7ql7npNxCLtZ
PGrbA32IsaZiJUZlF3M3rx3ImboGWVYXd50QgrGjguCBPj0UM1k7pg5DasFrpXJTarifROLM2ntt
UGS84UwOGd3/gwpZC59Zz5ea22tsrGyLldxN3oE3qCUZI6TE0hc0nq4Bn3c9YGRo7791yDOEyC0/
kZ6wIR3NPZZ9Gxj77ujhK78IXuEnm7KEIdJrxtnldP45xWNK45qDSC3YiXAGWqXRiR8EEx4CVGop
8lahfp2glyj1Nys+hOjdGoYS8cCviUNRVjz5Yc5M/WdydM5N2pYRLozgGnKSPIl+gHJSsdtzhYrm
jY27iurV47FBPbD7g4xp9wwiF1GJ3HfBkADZCfntdl1PiLODzSwRycoCitxtjzvL30TP1141yZCC
jw3f3XOZnCINHWL35VRyeDbVPajDYiMLZK3JgZX+HcVCjfdQMBd2mlDZThgj3uLbtuFXJE9T1rd/
oLvKRMS5SdxmReJdMs4DeI6hVx8DEqN9VV/HFoBZ5uRaKSyGBOJXFoLgaVqxdluIDuHNx0MGWAkh
Aw26R3+dwebv4Q6VqVinAYTy8KOB0Z7k6D8by3PqHNs6ze4aHevFmbK/5y2qtvarHFlQvSGvsF7X
yCTdirO24+SrXR7PRvX+hcO+VvQBeiu4GE9+iAkeIheJIEQ7N/Vj6kzuIM+tJ0XmZxENYevh62OD
78pdmMfYLNr2weDVfz8JdVQRVHcZ//fNn6vRBKlHOAZEG4BUtZBoLPfbjlVt/Y9h+FnHH2HYOthb
vG1JSLrWiQDrioItojDjSUc01vWYLKxgFLMt7KRB+cIw6JumYEib3VuHylmWLoVqWbHtQ9c/jIb2
/KtaA9oVAzFrELRcR7+JihCfjs69jOHfy5p8pfMtm1cm9KGWCazn1Z/wtAFQazbdZw8ChTs3n1yg
Voxom+tBvIXYj3khfLIJVfTr271z74nvI6c90Mo2GCx/6PyzMyI4gy+56Uu2ytKxS0p87ddU1pp+
RSrWoraLObjlnbEDh7TAlDubIgUpymOS3YaZbA6fKnTv7TVbGMxjVHdS48rsA5Zv7801OfjkTQFn
gqVHgXtFQOZ073hs6wOfDP9CdMDQYEtzvezp+B2RGhMkqXk57Wao3DhLRxoNQczSQoYxsvDIY5Mv
K9SVVb53QBzDGqaMoXkTakBUOYZdV7q4iLLyR+AnC5GGvHG0ZE1P6oBtCYq+uM1nnXc/DZsz5PC9
MnWMRFqti5Bs9sT6wQ8ySSBqzM7jfI8SDHxlfTTq01ZaKwt9d7rfidX8nq7l5gzl+HLvFBItcMyy
GvZhuYEiDqP8cpiR7L0rOXAMh1KoV4sRXvFkBwI3FAK9ZOccu+RU2Fpc1rbPc9P4xW2MpkN0ze4O
clCnMNueDvHQNNAgv3CywokCb43KkBcHKLx9FUFoy4O1TnP/kHd4XSjA/wXzq6EoPhM5Hmn2ytEK
AIQBpAJxjmPw0R8Nhm+qwID/VEVOrUUzCWZCPww3WGmuI8bj3RHQNsQIF5bEvIS/T+slX+fVBee4
GpF9VysXw1SxATCmlLs3gVdvFmx0kpeFM1iIg0NU1tRgcnm8c7McYsmp53N1vN2cJItN2CYW1f3/
wHBgfo3he3GhQxI8PvIfsrlETxtqDKclTAUcs82DlrntDyRhGEmFQTZSeZLlUOSGB8CEaSy0hkqG
izdzGwqiDKy8Vhui/ARdwSk3GsyKIfDxU6AONuN46ldMtuDKnKkZqLEun3Arsr+xJ0W6VcPtNAYL
89iSv1O1apD7ueRfZRbqjTCNfLXM933DYFKEoV/p6lGSPSrkqjzcfJ764USfCV6zGAzXcmdlWAm2
sTOpnnC0H64HR3ugbgdj9tiUU1GrUI/u9TIwqd1oZBYac7O/2P/qMWb609fcnMcxTF3sMce4xO3J
hY2tzXBlI9zjSsnjlWaXhuTUkPn/q57fviuZYyW4ML+O/SZTrhDapG5X7c6gxvQUdycktDw+iBml
6VUwYXlTKgL/FMVonaYwHH9InNoWGk4aN7wuTxeBYZt3Hr84Tj40ESVA3A7PzhOSsKnCau6DiwGv
yaoREH7S1rZMebk/XP/hOh8Ryd+x+bK7g3ZR9SP5dqigZq8thKD0/4U+bwybbMZO+yXVs+MiT9cB
7izZ3n8VhdtBjB1qBFaefUUne07K2C32M8MICGEQ2ixu9pRG+Tn+t5Fg1o8m9hkMTCh7i3eBrnNP
ufWJ4fYuNwmAFZhPzS8sBm1AlnmyXC67dSl7hWKE68iYkZVMwV+LC5p3J4JYuPA4rTiF4Rr9hgAl
p2IC65O14jHx0CnDw/k9sfPvxVVAatALDxC6iWNTSuJ8xKV5lp4tkpdrAQWltx2X9lfPQ81ErIRJ
Ujz/IP3T+agjvD9ibeve2UJonKd+TTDJv6K99LA0/yInoA87DYcPqDwza/InQVUUZiVxT50ziT01
QsZgSQ/8i2hz+LuFrsimU6G2zOGE0cEKbW8KPMy3sptKTcQNarMzpXVsERst2+Hf3NVJEsykd4tr
johES4Zj5QJH6f3GYfIMSEEyjYNOftVqW8/LuLNWoJGvT747lPNs+SdtPYW9VXxSvOrLPqgDzbfI
jtQ3L1FQi9NQN/kxyGLU8mDxHodnNANxt2yeYk/q40UutcXDvidcLrbdMawRfjBpUe0ZDyGOa/vW
J/7Pgq3deR82IIiUh1x5IYc58BADjFI/3gOsMdEpowpkXzIxR9vp4WUYfYxWL/PYh5iFVniRmttO
GV4y4dDPIxuUHyP1hlgFmJhSd+qA3b8uw4T2oYO9ooSDjEzEBsgZYrvlilAX8lYPm2iH0vaW+3ed
ebBoXjQXZQYt/v8PTcNbh/hC6bsah+D8OUJZRZAQ1Z2Avqr7asRM0wAY4R9qrgaVMVGZhKDdhp/6
tsN7heVSmCUWDpEWeuKH7iBtF/a3cGYoxHXKQMb8pNKDVy16CeL7w+riGxdlWXDln7KVF3p3G2gF
IsBUhWAj4LHLPV1695HZSc0iXgxs9/bUe5Emg2oJJV1gIkxvR1wayASZg88MEHiCQ5YiiM1/GpKO
35k1xr++dBQVzCu8wWCBobdyWLxNRS05DExVaCioYX8jLWkq0U7/DQmAZaqvEyjyfXtZNp7G3IS5
rzFKHFsRmBWALgn03to/Jd5646EE1J22kq0KHxPvfVRlfq31c8xHh8y0TW1LN57Pg6t/mCNFlcPr
FcS7M9lNUVbTmrJSMNKpOlXe3Mdxd3awfADMwcXQ7P7vEAyidesCJOM9hIM1ic40enyR3NhD1wQF
s9dnZchUpdDGO//juk4KNYZAxfIa5tVYvM39QmxdIb3TfScmRnqjCwhy3yNd94uXKZUMThp9CSYw
zEcECLr2t6wDpeZ2nb8jyFGmlUApn5FiQcVB5fUGljwqo3VYRbL+IKba3C11vAMCAheC5WQPW9ro
7QCTecSbNepNMM3w1+9pnatvJ8xNqhunEMkWdjOYJNZWYiqZDju+xEs3Qpt21uZ19zH7zmdQGqwz
2LubrWMa/mtF4xPbP4sA2yzdkdcboIBLj7qloxMAAf+5evzVc0uBYS9oW5nOOPb8wWUmcWRkRpnZ
hfw8zFLTZ8izG3D9oH5GfArGHIflXn0zIdjBSZEoZzHg1AMEXgeC2bRZ/kg7jo2ba1NqPt40XRQ8
AFQd9C2VXlUS81jJHwBgnQwLH3g+olSBoUHcKAT9IWrHjt1ITeAZiaNRe1SkBMUNd2ac+XUZ8HKn
D4hr/zib6/haRbvlZKtP5tJ+hm0ZAPQ+92lrdv2xdiJ7Z3zbUAhS4a+rggQi4Pf3v1ijsQRnycJu
xpqKoE7Wk/5+1AdVXDgmnCSuA9bY01eR/Y7IwKzHsRQq0D2ukzMWM/T6u2Dw8q/7QdEGke0w515O
00E3DuRdYTIXFN5IeK7vMDhS0t3Fsk1aLNQpPcWzwfr8nyMrwmbxPfEJRvcvXWLboNxPeh20Q6XX
kVwJZfn+u7hNvB6jKRh+4flBNgvZOhRHWWAmalss1xOaUEv4dXiEBI7s4JEk15Lctp2XvfXVGeP3
zT/iYshmErADpII6Oq8/njKIEq5QwOFifXs9AwNETPu+JN2J1Kk1ptd+Fuu6ADnMtB/kumaYvam/
Q93/sbjMZWhyP99vHo5Z77iyb+H2csRsH3RjdQVuOgOOHZFYQ6wWuDNgHC3zDoNuuz6d2gtyJa7f
3TaDGUaIq9R4zcA8UjnTeWfcIw+RKA9UJn62HE8APSJtwFYkyaxAKzLcbGU/Lbu27V6Hv1s8kVRt
TfSyjanfKj6QyRRgsRPAg1Jb34z+6CjmowwgfFXXWKPG55O4AdFRLQ00IgVwe9PQ4dULLXlc1rI/
Krd5JNKpcvX39eMIkQIJQzUQlT4EXiQruQEUMTdaRLhbyI6RtYj7FquDu2eDarOdOIA6C9JbAc+U
lcXZTSHOsbu/Zy+YJm5aKu+S3kOib+FTGNY17t9qezc3HGbDn+K6bHl7lbrW8lZesUR9nuv9fG4V
v0IBgIgfpDaI+JwiOf+n+hHWqSPe1gbZVmUTBZrkNH7K6n68Vsh38GrcvbNgZJoopaKxCbijTvVX
TGBFaDVzA4OO9Du7LrTbjAHypDRLgyFuAWNtwltsVdyp8F30qkPYS1MHqS/idnaXniXvCEhJPw8C
GbWMcruDiT+B4JF14mySGxeqvqHCuPzcX6+HSqzUy3az/BI+tb7uumwhpTSM04vQgGVbdeSvErZc
PhFzqhF+C7v2xadce0Pm/0ldaeKe5y8lL8cTGqlXA3dFmQ9Mbp57AxkMXTNbS214FGXpIf4r310Q
uqTMFW8rY3oNn3+jxQ2UMJgLm3e29TsBhge12e8dTZQvKIoszyEsww02yrLMxiHZjhbYKaNa9wqh
8EgrHYEP3P+g8l+Bf3SfL+FWOwUbkxT/gNLYJmivelDHjxbw+qvRmdyXXvr96riJ9SKjxdpluzP9
L2tBsMQYMWl5/2AxzAzYo6ptblv2ugyXnLbFpqrY9LepFRQbz692JO3xU9t6sQk80WouKNW1U83s
SZfRW0RgV2BjTdcIOHQq3Mn7nNAdZ90kvXZS4U7KGXKeFDGRmb1DLRTEITDhe46/ytSG3wVAD22o
YTWpFwuMkjfRq8d0Cm6+G80zynDAv4ulXNEr8nrFMLItFM2nC8vsxRRNReNQEw/MiIPIUg/BlNtY
SjmM1/S5CG/AhntFHSyIC9KC1wMi0zvnigBIB0A4I43wGuZzEttCtKGAUbcEmSplZMofg6hPDfZQ
mvVx56oC6w+trOlBSyZF73iCIxVhivy9qOq1+AJOhdOVNGvhqrDAEq9bcrU2DUZX1QaeTaFGnpqU
VedKpE/RhFxnfM2jd+FFjWTDaOeO1U6JIy2lkGUW781Zq14tWNqbSvZp8ZA6xDOePPQMcEqtykTV
0tstrrmWLe3g6usUFKTBSw8AxV51T2nIKIt8xOaPIGg2+H/Iy6QVoQarJTUw16RhblJMXSABcKn8
ArTRHQR0/TsiOyBG1AAyjq6/zsO8YXEqzXE1UrJchlxGbliIyGvRF2upsU+TUnz/NUrB032BVI0K
emnhL3pdaEM0hwB0+JwIH7kgq33xBT0/lsEAWaeBdldnjdQT6NehYFMTj/UgIt/GYbeGksLp5ZGO
tMOpbwJzYmGwUM5TTb1Cd5YfaPUCt1+it+gibsRdP5hEHEyk/9BSoUmBjCUZjYwrAwPy/tJTzfXv
oTrASCfEpAE23cJRl5ZszENDg/qpkx7xpMe+ClhlSvqeQgE+YTNTfQwRr4dGNlIevD5zAQj6Dr/c
MSPZzWDA6hVZ/RVGZ83d/z9HiZ6AXXH8kTlPonLtLfdAzyayPH3brk4i8nE6rqBiqZ5IJmVzroZq
wyrT9JueMPpb05xJyhumZohVPUGRSLXIRR+BItgvaLDphaMja12ncVAB0parPofgKJzkHKvl98A+
D2SYYMPqav3KuAHUvy4hsHhQZSwJhwXk7eVajOFlAls4VHoxJVUbTJJy5maqhZImaZUERIcU4vg9
tjvfRwit6pfjfLqZdcLlHCCmIQdkx03jPBB0pPFDdHQ+7QKQ96KXbAh+PbJ4MI/gWtPTc+Zbv7dD
XVi5ykvfCKni2mlJPF8YcDM+DIbamzNH4BNhFbGo7KD+prLYyiEwJxXVsBLF3yTZilV8kC6MNaOh
v7dxf/UJ4o3F0HVnlFbOkPti9LQFWVyYjf5pN995XBVomxk0gFH7aROi/3Dh3eOvS7z5GIbUjGgp
TCR2TyR5xv+Wsex6g9OqgDGL/YK95xe97OtZhGdBIwaJxw7cMN+z04JIhicVmEL0rT4VVM8y3aWh
JxYB4zVmqtkNWtyK/SiQdZip1zMLcwnX+9UM6D688k2AfLqiHFLnvvwihqNbuOOzj8X8G4aNmZRE
sRQbK0C7GQaNmLBRH4MFmF4kVvIrMsfnO/AF7OuMMpmAc7FXSLLuCykgtGp4G7faPC0VZfxtgdsl
uJmbtPrgFw9jgoQiHt9NuITvc5ojA2NAImgl2III45ktE2uiCr6ZROR9c+BLx7DNYdekR9P4364c
m+YIJ++IcUGp3L3wKLBjcjVf2EXjMuJvw/DeUhe101yxv//JvS56XEvWjfBL3aH2y4/gAuu2KwQI
PfZOgkBjylbcjmJdwcjKA9ktDbeqs6rnz3PLhEgcL9x//aUn2JaBNVZJMcY/9NM8NYF9VoC1kfLf
IXCjM/ESigh7p6Y6yyzuQQsBUyx/a/d/LfJLFj2ewW5COsLTN7PFypZfQgjEUeX+9mFoNJtV9UEz
Zux9QB+Tr6WNMwzAEJTMDpTzt9VFuqLM4DvsoCh1TuKjjaTaCTMYJMcOBMpnbsw8wGm41745CXla
KOokoSGSJZHXt04kTCF83gceObjyItgTz2kGMtCDJoGxYtlKT5lCuJPVuvS017p9lXPfmkyaKwFb
r3/6KR4v+bxbtlkQVEjKifrb0Cb91HdWWPvsC8jKBfXKTSzWHmaxH7Q8TAdPNr7D5FgPViJMZn91
8JcpdjmpJIiKAAkjesQ8hjy3U+RHncNb9xyfu2xf/AMbTIxfoA2aUWOkqcI6Gcp7BW+1T9qezJNL
wJqYf+fPknITMcXijwAIk8L6awkxcNXKyRooWgtll7kuztSU+ELqjxiade/joib3W+nzNJW0sbgu
PSMfgLx8aFO1emaM9T89s/vcw5edze71/wv9juQ4VWOTdwOHwuB9G/eRhbfhubfvK9MZW/WiFKhU
MH66lk8uCxScBRsizyfRC0HIHYOhiFx3tTmw2pBRf/MvkQtKHaVsgbhXkj1N+f+4JnaMWFkj8tnp
46dk1BckOAlE5iCl3y4901SIIE0HDV/B8S4w2lAQgHE1JOUAV32NE3c4CGMCuebEJLFC6tES9Nfg
xV8BxKfwuL4dfnQsrCyAXm8pqA5aYqWI8JYeqJhc9U52Yy+XFVZ23uUv9zxqvP9t/lNcku88g43G
TAPSwzBGnGVnSLMsWnI+3SwY64xFsJ11NS2MCHQI/kCtumNt/aUqqYa1M/tyFybncz7CyZ2UrV2R
tUyFhJvmNGnLo1PMw/m6RL3YUF1uD3O71XlJUimx1Cz6ZZT8OEzwqFvtF1vMs4bRYsl/UbtY4Tq4
KZNq1a2zozPglEloIySaEj4gX7sw8VEtq+bvoyhnza30HYZVfzk0VM0O3748w3vi0vlxnL3oH0cm
svLOxvsvR6rclQywVNsf1LywT/kaJSIeo7YbgJDCRJgTxQN7nsqJOxTEpbYNtbiQ6QW1P/cl/LmE
RGcqFHWzWGP5S1YBPRO7XYyYpfc2rnb9PTY68JVsR2sV1Q/CPqgEZeZhZxEkoAMh6XWCMzUH8/Su
LxSJtjiaLdNLG8k4hmDjYxCJm1HJ3lOmY4GB6AwUcwUCtKhS1nYqq1z0DVPWciTe9RmdvKUDpOh9
JBDcdeA4A4tTKHxlLbFlbmdSCNa6tR0zT+5eYrjjqhpKXNKQQfXNiFhlB2jPI1JlOG3w3sU0LPet
9raIVf6uNRsqgWP6cGPxw6PvPHZsyKaohcR6ubk083W/gczIm43yhknZVNI4G0YjZbqtYRSLHzwF
Jbro+MJSFjzeCvo0BHBY2KGVrAzJZj7PWaTRRJ+nsoerW1ZSjQlvMHB7S86tFFqlqljJAENMYM/V
PJn/5EM1jKq5w9JFf0hPQsEzEPl2SEkHExw5Z9AR7fdEbnb71lb3GpigbFNk5o8O+xnlpkjsGyUV
EdDeOTBGU4DOkHcXbJ9QaWzVMAhE9Bn65r1dQ1xJ5yquVGc8o+ORu4U1ZHcZUHiyC71gugaKluKy
rr7b82X1byaPwpCNnBem3atfdLrP/5DXT1PJW7wi3fUMeg5eYjLzIrmI9vI9SQmK5O+yBMWZtVjI
sRvel3fkop9w/z8XLJSSayn32qO1FjBOELzH3kzJIUKbRfPUSZ3rEnJw
`protect end_protected

