

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HZg7J1eicTLULECaPz6ctaw8y1kpWgApgtfn3Q+zYY0GMZZHrstjvvtt0rjShEIyHEmHswkTon9F
uInqopAFVg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L2/HzTdtpI+DDWwQZLtw6a20VAniDvlrZ5k0iYB4G3h22Zth0ONh9GaVxdnh5RvsADtDStl24FLn
89acqSnMq2//5lAdWAp/jsSUiUTqUuq3s51XcviRecb87oOU+8iTczHYM6EqTAd3Utr3aKQ7HiMo
3WL0mQVpCBOpCQUD6jI=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OUJeS1bwtebGQThLvBFH3PwBsgx/p0nU2VJ+e9SC+Hrio/pbJwz4o2xpS2Z63xJ7QN7VhCBN12gu
ZFY5Ng2Sgl6wTkLeA9Vhfi5uJY35hY1D9sWB0j7MhUUJxRIFWIWs+H/FElpBvWn/H5UtcrDSuhP2
nLymA6ruYrGfx7a8Iq4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AkdqgHhBI+1kEGsbiaO9eH2SWpUOBQkGBwaPxgDJYtBsJdOF2T3rxHzMH8aRRo4rOV4wq7F5qDYZ
2bRKyZlKyXwxOIrgHQ/aFSyCdbfrrJedXNOvayf3bMLKWGvmkeKTZFG4ie8bYq1NlzxjEK5tXh5u
do6EoDDl64fqmvjtPSKx4xrYKjkfDGC1J+lF3Ws5x3iNXrNkIqRirBHfL2nwSIIbCGtaZ+SRJZcG
6fOBaI5sglgjVMndkM1UDvQGQg1m7SekmV1gNbuTjfVG4yDcoHwJCq9TChQTCfG05c2xR2kyrVm4
vPlYfKMD9L7sptBiihT7k+285Lhb3gyxkn+LZA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kU/KxTFv88aIggtPFaqaw71mguuPJV+CvKI8SqHLyiEfFwnEl2rRaQjfKPPKVY+a9ar3+m1VrJZq
XyAytb5FrHwHwKJ8PWa7bc9KeMqYCg0WQyqVAR20oTRysvr0JW9ZU5xcZQIfn1WQOAidCGjGERXk
D8J1Mok2babDuVuQ1k1BLyAGty6ATMVk3dUAR5LIplcmY2dcgXHhvtTjcDGgu02ufeeeQgDtYdEr
XxPaZ/IuZu3RKlqS+LyaN7GLtQ1sl1FVJL4oxiYEefZ24cov5R/2KmrDI47bvcitqcxarcKhbIwt
EegxbadS43xqD9JDNFUAaaCu542z6SRuS0zC4g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k6DApHKykfoAVe03+cLJSaTvIyV2mgyg0ee9r8sDTCqvO5kwFuomMl0B0cjUO/4j7+8GeD0YVUGW
M2t6DJMbIxuNlNctJRXzSjxwlBu2lOTLqWCd5V9OOHutCH8JEU8ndSXTE8ecj8B3ICDoE/uYntN5
p9eeS5YN3Awwuuf7vpsiQrcsy5iqvO8GW2b0InrBhe5m2bb+CK00dsnS6RTA0bU4RH+b9zcISWyN
JJFEeDryWX5A5kyBX+Em8sHpW9ssoOlBZUuAR6sGhqbdC9endcp3vkYasFpW89RPhQcAE2DOJVLu
qXK6y8bpxJSgUq7bdln2TJUwnHb0mgJEbAKlHg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 114672)
`protect data_block
rVE5YALEL9UfeqL5CanomekQP8u/BHYBmNdEWMt6CGbZzAiFYt66wyybX6jsrtSuIqPHUjuqJbPA
TEu9u75k8sWuDJEPT5BIk+3NS1vXh/AmYTrtqMMgZJ7k1MBAIoTW7LlphRraCZxxyYfiKcLe03mA
TWiIt/C1nvT9UZco02zaxxoKlLggP87jTxjRZ6y5wSX61uW6C/yHb99a3LDMxYx02XwaIAePkkBV
BD7WxZ7R+I5GlvKgMNmYnHxGJhbsddbIcC60LQS0tLBGUyHoBKhZf+PBF3GuUsgN82lVyyLUUUlJ
CZ70FMfYJHKbrq2x97AQi+z1zbJ3YPIO5N/DMaoI6MmR3LmSDUYU16A0lTzT6qoTphz9KvpGr64w
CtCY2zlFEk70vvWptkJ+ip1qpUJkmLOQndX3X1RwPYvmy2fRmI93ZQj2oCXFcKAvt1ho3sNU1Gzq
xsaMroG+gysYdRQKGtRf2304NKSxVhRfIaWnGl30SPxKFmCEWP8yzQ0mskauMQm/qe6zZPkRDBJi
wlAuzTB+9LQS+IR3WF1FT2TnfwcT2c0h9b2jD9aS2T2BdkhJkAIOGn08pcvB2k5H4/8BMrdxq+jQ
UYFtNPY1BQLI1pAR2JVu9PHz/Qy0vnIThr22qbCGszbNSsEfT3yRuT20gfcnLhIW42VWEg7YJOmA
SuxBRR60dZUIpYmkvE/eXlDpsI92z5xYHe5tQ2HdYR0xye87cZhFy/2AwMHwtMlGIIHRyLgvUIhE
WfEf6qpepQqROc4D/ba9NytJZNjdjvEkTtGfLIbua8QTNF7Wwp3Z57VG1veydNIYGNaPXJtp/6xA
CmZZqFWhdB5yHr4e3T192E2iAfXMQ/c0SaTrZjpJkWX0FeuslzWx6pgJ27Erw8P6s5wCCKSurhg8
GdpHT9PPhKk4HKd7gl5jhnwJhE+1guZVMkt8CfqNogcvYyrtCgEaLhnC5/+pXhZ/m7eGfTs6OkRI
FerAYIg9bNVgHqjhDaTQD02LMETr0en5p7HWdSDyzWtw+qucgpJ0e3OPFOMWUQB5XXuvSIjvlK4X
5Vo7+F3jhLfw293MVY5tX8Xf2RwwWguuPnGkotsnrNHqI9WMTjDC/wMHdTqMsAyk+0Fm1CVWSUbq
NS27nOIyGyATO0Ft6KnCGEUfhOxVItnHnC4C3f5H1w9MCgOxRS1Rf6VKc66bA7TKbmCYGosDKz9z
gPFr62DIo2rPI3pK1xPw5I2ULPBgtx27SLpKemeqBtSnc+t/sRk4uSbJoDQ5eC/KEynFSb7ThEeV
ro5pzstOV4SA7vn0znfDSLKN+qbfvBfm9aDHMeCcCL+b4LplEIde3N2cVT2WCAYBhUfBSvD5t62n
GRT2hSlKAPSrFPC3y6yfu2QgcisapTd4uFi3v4T3SUVGarHbjtxZkfkv4/ksACbi67yzwn8dW6y/
pIzNG8V05meMdGfOSb0LeA+gApHtkMrK7jNEz94TBaWdwDH6ie+3/r+6RBVzDUU6uNAq3dtw6XHj
DPmhOBZytECp1w9o+Nrupt65amS1iwXJIwhRF2SdXelojKfUY8M9WJut+Msu9+A3JHHXdRtUikMs
6ha/KMfVF1ssYY6lQZBTD89X5Wu3BdmDrtwJ9pvRrH5K9sIkgsK6wduktrPceLvUckr8szNiHHkL
BDWbkrUN4MB/7FPlTBzXmFxC8xM7vUzQAvTdHz3/fXP3VSoqzVfTgDJEpUq6/IpTTvE6m28VBaZF
lQr11ghtJZZ0gYY/hspnMEGZpYRejR1EC/HPgocDmS7r50vPk3kGl8fis7nPsgQ9AWYUxEBPcqZ0
UdFDzbhTUzoHI1ykt7UrQtEIMxgcV9gDx5ocZ8ml2zeqDJUrUXf1ZcKIgFjf5SmZJM7dMCxnVUEM
qYm5wQXHobm5sqM4NVwmyBBzIwXXCsln9vPL5J7PuZB5VyaVAGk8yrmk7ubd4Bel56AAiG4X+QLh
XtsKXOCdzFw/XOdW/8aVkBa9IE8ykFRQ75qm7wbwjZPOOnct6tRNNWze7NmPMUByCeh2PJJxlFKU
YZw09HBvPHw+ToLQxo3JIYErVau6Bm6G6tNWpwBtKLacYen5kQD5n0sF0TlT1T5O1nMDEO9u+Xze
bgvt0grFsiJnD6CUGZ5oTFKGbN8AxKe+bZKJjBlKYlqhHZ/3C5xJV4tY3P5J6mJPlY9+wnEvEFLM
Xp+ZGxNvIdf/FTg1uiWv2tbDLZ+3Cw0DUqR1OeXWTxh556iMt1i0uIIx79+ChXYviJuA7yWVX0bi
KYAqSoBtg0GrbCL6f8fzjXkfGGN8TwN0WIYRuWh0JhHC55OtRWkosq4d6Sw9ExIPx+1WaM0/okoZ
DkBKaMATTwZImwKGJ3oXrERfIfjB+dJp9E7frm/CXZtfTfoUy7lo8LRJ0FUK7wn+b0NASSEYw7Ug
Hix/V2yY8Hg9AVFjo6XULdzmkxzsrKo/qdGl3rn4qzmGNlXe0SVHwvQtEFTVSSBttIJYpuy8L0kY
iqVTP7Em9ORHsyDY9If4UWCY6gVH5uZHhDeVl7WTNZM1lz+Ph2t4YcYy2DYFswEFdH+ot4pyZ3CK
yqHy0Z5KrGiEsn/UYF1D3/BBbU72T2rys7ExvsXr4EoYdDCQgZRvDkGaGj0/3lIWKex0lqasnDQK
jf1PWvT/+zE0Zv1/dQfcgdUGxlhUX81uCrw/Cqi17rAAzDPhvTL5/6EsSorT4OzIy/i3PleLszlV
JHUzZcHZa1N2zHjBhl2nzgnnpNsRgeOSynf5cZ/9WcGsKvLgpeo4vHbh3HOUyrFvD4OYe6MRA0Al
MOmbYPlGy1/okF16DGdj5lDofLLl957kyLBp5ccMC9ini+vNf4Doq7+VLDGn3zY1YxZLrafpsvnJ
K66WV1YKBHfZe3stxxceRyRcLonqzLd4yoXrhdk+Si7EohXNVg/hA7qrF2F1I2JpflguNfl8kpCU
n5xO2rqlCXeTv4eMP31iN1ON6CVrUI+5BRqoL+NZ1+pzTJV1JaGjUASmeh7juvsxVEfnRNaG/WnM
6kwFt6hXR90nm9n10Z1Eg8UnfnW1Qy4owpGKeVjKuXOYvV5+vkqJ/ScJTSwpGvVt+vdUUc4i9bt6
h6whPwbYHGFUwR6HZG+rrhrRianVLlzj0S2gQwZeTIpDezt8yCUmYWd0WpsoqUx5NiyxGwRiGLCY
JjmEsWA8tIOW1VBsWvAZAp/3f9L/jRCIQ8nPZ7vJ+obSLLAFnL6o0O9ZsyFDVXOBL8O8WpqLCUQp
EdJt7eWhoDngf9FIEWl1IE1z6nFkNZCZHQlUTgek14Q/5E7uh3qeKXmfi6Ug7FcE1hpvjrRYVMAW
EcchPdoc1DJjRwBqmMsIMud/mTYNSZu5YtZr9vDSBCTq+6vzMxSXTEyPvixDHq39V/c/kGjZ0Ai5
pkXqZwSzLQgjRr9j9mZ8DSecQv5d/ahhRjA+dlsEAoA57FNATjUdT+IoP/154wt8iSALUWOwvpMC
fukXVRKkoFr00K5qjlVisjjn7jiFm33WJ9HWPsC2CVCNg4SfZVQst54JA9MnDGbtpqiqC0G0K+0X
kpjvDojdBlIWxWx60bYCbBc/CUygT/+3z6TlDCO34cfRR0sZnvyJluHIscnq/Ohm1SBkTMKvohHw
NRZqwlzvaIT/Tjmluz4nNndrsmq6Te7wQC9+L2MULOw3mdaiHbiF2dTPL1fdURmc9xFOOWgAXxir
qt5x7UgqcYcVdWxQED3LHQEZeCBhtE70xBBeBTojqM94XgGw5LrHcP8pmJorvMpRT3v3GrqPKUtJ
YOf3S4z9Wrz0Xj93qpuEWZ7pedAIOXPlHPBpcbYwlf8WNKfUie+j451Jo5GbMFHnAL3Q27PNnRCl
LvWuCXWlzX3J1FIGNjkf9WHE74NSPTG5Kb19yX8V5KZD84jY1jj/CRkNjKi63oyLNWNZTY3GEXhY
h/KDeL9JdT+MtyLy4n4qMqMjv1O8epMtMcALRyIWwmNIAQSSpTXJmPn1dV47FD6JkgUs3sKmReo+
VwZXBI1lp04MEWbeQ5IJeQ/L5tT1Qd3nNQrY3HefD0awHhURy5+74yk4lpkJqpPXZhPIxc5RpFyp
Vv5WKpGlf6sfrlieNlogqq1joBNa8ZeDbDHev9lDINvUipHaHDkhrCHYrdzRTreFTAQCf1hQuf+f
ruIf0MIPpHYEdZ4nfm3s0AqtAf4VaK4uEbilzWW10HfFUaqaG7uo75rRdBtFaXM0U5m87ki5EbGi
Ellzs+k5eKppCcv9SKrMxGUOxoEiOvUr1zmEDXg2TGyNR8R5I5PZDecYMKmctNwY4zo75xvh2hPH
bgT2quByzt/3YK5Bk4kP3r7/5cV873sqysk86dvHDX/d0pVfyo+2aWhNNqZaqiCUv8yLZ/a0bLLJ
MHtEBP2OUZXCKdm+2vU+ymHPReGDBYSuABOu9hJsgjaAc9YDmVzD8SJCry3L6cqWHzcdDyN20hfb
2lBdCloeF72tEOQ1qrgaTFBw6h8a9pKbExTHAFk1QcKpnEXR9JQLugF/6NHJG6tzWo4b3oZHQ0Ly
Vp3fwSgeNzKpmZEKhi98z2H/zrIF+Q1cCAeuuV7ZG8nUI5PLPLpSqYiF6onJ0XPZeatNjncAjy31
DcOEia0XkeaayahE0q4THNO0+OkblyYeQpMk80T1wQU1iCYAMl2dX52TSTdNYOL1LcTKoH6hPivd
mmIJnAplfOHSFdLp9mTJGD0ljZrxK/3c9rV9Jv4Vrz22oxmtu8ndCs9DqNt505TiM3KLcR6bb1aj
5qi7hutrcNQx7YUj3P/2CtJVmwyjUJ+Eejx822LnRSplDzRvQIAo7LB43V2w7/6eiRz0+jp6bofO
8hC0CNUdXls5KRJb65PgYo1GsYQmyGi6jdR0FzT+pEKmLmQzD/16O42erF2lqVAl7wVFpnG4JkD4
4ml32fr7p1Zpzus1xgUXqvgtnIGyPvxARfZma03cjjiLEwcz5w2TJlACTohnihS6R/wfhaHJhf8W
qzSWWmSeib1HjnTGH/C9rrBjrbrJYSebYhH+/xU0AoHRpiYRPYO4/s+6v2V83mk5bUCZXjtrIBsg
ln/6MNer5EORNp41vPGd18PwFW9KShBsF5Sv77NOpXljbmrmmPRfgw0RtNzfszgPXDOs/ofvEIuW
X1eu06iw6QFHy+1RkAGeDBqUtg4WJ9to8Phlllr5WK2ypTIhuL8VI9NcunvBulQ1nAql3D+MRj4O
5lPkJnKMMn6aNpliMAgBEBvUEs4Fv7ZSK0wCB3Ldg7Wonk4mK6NEV004rL348Qzih5txjRgLdubr
hrI45xTJrnKjrr/ojnGhTqwSeNEAGqtXF6OuWnijkPBCzCc4h5xWpxSXtDgzMaxDLLsGi435OiuQ
0Ej4vXqs2Bf1xU/43VrDHQdHYAXns/ZNSafoEME4ra9Ze+ke+MlHzqZquhpcLfflrPp/OGQhcFdr
117Y0GBNnJ3z1JzuYHdJKz78O6wz1abc7QnRMnFPy0TpgQ1gH6M0b/pwKnkC+vJ8+oOoNAFXRdTT
PPtcWpkD6V41p/n5JwNf3ur6Ai3rnjsPaJdtJ8l1yVL7WLbXZY3s9sdDeODIKuc0rmoWwAR4JDnf
SklUsbG3d/7p7Tfug7p2rBuBhkPsCT9pZyMggmIRR4H6pa/Yd5r+lkFx0b87tufto3eaFKVCPq4c
GMCXRpRX6/qldkWf65TvwZCpHmjRq+Ojc9yDa3g2+hsBYudpdqVBmR3CxknYTmcZ9DPbMYrQVRFv
8P/dvzN+BHyu9CeYNp7WPPpFDNt+sbG12l1G8hH/2JbV7KV6azw1cYED/czLsdzk910Xh6tDNerF
sjm8zXxTa8Fd8WeHT53LOT/iF1rGOJ4Tsli8CztRPmftrj3LC5rTW0NsAi9DvyR7zT7x0Ie6mWRx
gKHm1omfvFXKUOdk6hE4YNUUZt4lj6eWcua+R0ZIRC42CWiuXWWN85ab0gHDkZH1jkvhzrnTrjqB
PrSzD2n96EUzOxocrEmUWwDZrNNUcLB4/Ua6OUYa1Mju2nvTvaZXZwugOwb9pOs+OEYYCMVErvDc
i6NiEf8BeoaUucxjjk51xHg/FVkqLiHjdaa9TR2oJar1txeh7tEL6XCqQUL52Azcsf9x78fB26dh
+val+gHvWnPzQHKty+AATGRaTnXQT9s/7scNBTWKKIF5DRTvi2AK8T+Cs9wTkm7PJ1MjFvDrlfba
Ai68ZxFViimQ8HfJ63vX3/bm3JpHXqSDsG8SPCpqa15gy6xCzSjVOARwLJ6qizdWouH+yDi4l5rD
Pi50S7gww5DiQF9crN3mGYAFHhal9maN1Y5XgRcgbrY/IJk1pPMl6HU/1Dc2Zi2BBVVxLylwhP/n
/TTcj8Wz1MfWef6gjBmIgv9Ly/O4+bUk66+D8/PL25GoLX+cTLg2VnKqD60dukwmFhXJsckLm2MK
q1JNhTgRaAwXd/7TXdpcjFLP+H9aSrXFK/wMCZnKSGwipbujlUCJ/YIo1mKIp4C2K5fJ5zLE8XPc
Hyy0WTNieU15ec0sfxtHIzMcu4tLMetl4L+/cZJQDf/2bIDOZDJVKJHcnbAV9aDoJmc3HRIzzPLh
Ykg5ywW7ezGVXcT2767426MsZrwwHXe+Qg03jT3dfuY7mIcLGSESypiF9DQ+ym/8jyrWs7FoGyK4
/E54MvaIoahG69voStODj6sQAcrk1gapHS1BKkyqoRRTHh6hFKQqnFMNsWUaO3eVnQTGFnLhVCLe
2A2MQATO53mjglX1nhE+U7gzQJ6PyD9Laiw5WBwo3rqLljXVm7sSJEjvyP5mCGXrisxyzFot7RGu
Zvst0WMAwcLaCezPqXKbM2YKfB2jo3AsTti70gWhRRznvT4mazSnaZFt4Jsxr3DsngbUHhisahAy
teWoGBgjvhkP+ptuUjxaM8sSIH3LCDgPzUgqksFuMj7S/e8KrwjyawuuUNG7K341hfSJ47X1arrl
TwNN5WkczS493rOy+6y9mrj3Bc1NsTdNslZr/UDiCvlrfJERTWBffiDxt6O4Vgb0+QtpNjAfNuJQ
bZ/OqJqIp6U+5szRIzq7aZ3ZF1SzBTh+9XpJZXlWU8KxQH4yV4/FjO2hjwPShmG8GOSlbuEmFztJ
Nt21bLbvt4z4OaNr1Fb/C6grSzbBm/LVvxz0/3Z68mbLbcoI65AyxUYWwPK1rjzm0XJk+2kB9lxg
yj+Mdg5igfVrRCH6fHRrudKfPrVSoARj1lm4yqRAv6p2WTouFAAD8oVlDq4rLGhV5vRWC7rpqsHW
yDtvqab6Xwe/J3GwOPgYeyOwMVjMfmDLzsNECxeKSI9fHiS9WEu80bgB/WNMze0bTpAq4H1oDNvd
1MMPtbujpQZIzZ+BEByo7QoClnUxqzSfQz1Iu00v6Hds64D+C02HiYEiAel4R4EB1f1Z3Rzobosb
aP8OVsd8aidqK/Nfopz54oEgkjvvK+i4/tcJrxyOgNe/32K48YUPev6jDmCUUUXXgPG0fKeCxud9
spSWDp/agx4duLY44QIJFT5rNtbAEzoGq/NpesZlOT9YS4TKdG7nIWK2yLxuyoDYjpB+Bthvk26C
b+subsjgBALHunBAcptROhR3D/izkl/qcG2bYNehiFTK0CUVtDowJ+B2bI+txUlwox0DH0VyTYrw
YQkHlY+crMb0ANqc+LadacVnvpF5evZhuZvcOW/PQankA5d0W8rwYc2Ar6yLMOLnkHgOfNuSWVip
KI+IHk64dYJnK26QosBEkcB9+eNWsJI1cw3HtHLvF1edrzBuBtgVXfi+OD+pCptW4Y7U91imkGZy
RptEw3DJTJ4yj6RCDA5yV1tSC+HXS6yC7GEla7vFPlltuTZWOAOJd9zhW6yYAPbTWnkEAxhwGm1d
nsYTntGOfto0Kab3WnGIhHpNQzneLvTzlK4rRqqVQlls6MkuM5OwF6ds1HpxTYHxjqfS9Js1q7K8
Y+yixdc+6/BpdgfanLYnxksgHNk9MYj+w65JrcDoRnz8iL5tIBZPig8Dpvo8QLopTGMQIREF89I/
1GErToBjYzQoj6m8rvFwuv7ynZ29oBeUyYQ0Y6gSyP3dYHZqMuq/i8ER53EuJhZu93lcmkJpbv5c
8P7QL9nLhH73vxQZcYlHMkaHzFV1/8NStdL4nw8xw2XcYsJiMXPlVtPhKnrmxjwjyhOOq9iLiP07
x8Qr3tB8mn/YW2/7cIHIaBFbNz7a6BCh/ys6YLZdquI+eXT74mu3+yy4ERDRhE+Vdpix/7BG/4m9
/gzwCl9M+nA4xU/QqKPoj7o0eyPsuZDD72Vx1AO64MTUCLcuH9KtldPqK73ngRBl1fwqd5J0MGK0
CTMhLy3+Hl6eiZRNhoTIF71d/uR7R0ft1J+fUL84GK3yea665e57DK+MupWWW2CNrwDFOQpbH0Nb
jY73f3GPKjkDxQpzhYsdE0j1cU7yQ9BGh1gcmc/lSqkClD2WQlKPa0CVKpZ86ICtF4oSl/9uYtXk
f50lf6F8yX92jJ5PlhMnZD4//WGMVI2Mtn+mu7zNi07LWcnSsoP+Q43CaTeoMriZAL/WVzZbNNoF
mI+f7fhhwDGcTwAs5cwey5n3HnP+MeCpuZgIcMDouDK4IElee/KiLenFvVJHSHd+axF7vRYudsRV
MNlyBife93bD/CTBr4gsRXRzFCjOhM54KkLBi+o1Eg/zaeZU/He4e3j5Id+LUKsiEVHvfeeHM8/0
LzMunoW8gSGVklr0sUMez/hOFcdQV8T8YV/uZBQK+rrkJB/MIhhKfufF8Pgcn67oUlfc9uOG4rze
M4L1ybbkvNutLA5hD4WVBU98xd7ibvRaaaiNgPex/c7XFgSoXIJ0DPwmOsE0DbVJVWOXBDguk2YM
JHiJfjYiWhJHjjaouuhsheEBIrspox+rxY84ugAM83UwOg1lawzSDFa39VkOKa1ndJg6OHNZ0N7A
JbKH/hJs/lqHR8PgrQkz6L97lDoizSy3dq+04EJWlECKKDPj3w+036pFKcQqzjt7wnZ3/uejtt+A
2wXWk/WiphVXlWJB9G/xrE7HhuBp8WwYl5TEGuCqwtZGQlpGijfzrv/KY4QWdzfT2WPghpXJauhO
wYez/dI5RRh/NwMmVocJuc50kJHnjHjXEnNQlJnZJJ/7uTNXWZps7M2lilWnNv1RAUZn8Wl6zy8N
6CIRZnRMajjQD0Vi0ulN5xd42lTgC/o0IO2yCdyn+u4MjX+ACxkkJRCbeoOO/JS04a2IWJYOMo+g
NUFaNPaGEpxOomvwWGm/YLZhajw8b0QbuS1O1q4FNvP7DpWMxvrC+OeUZQVVcb2IBKB+1CaQDDks
d92z+sQBGkC+iFSBN+vO1OZ4/JNE62wrEON9FpMp45BRNEB+AxzUSa3+rg+dScaZbWSlBPMQxvFt
YauG5YKLX3jre9g6cZTAwbfl32knh+vSHtk2Qogi+2XJejgPiSbSE09kna8nFpsoNs4X64SdKaA7
siLFgJr0QCL2KG03W1c0nZzVNUfnUBEb6Z2P5LYsC3xPA/i8Wfd9lOTvbxjoBaRyXU3zdipuc72W
KudetO1C/Em8LojWePqUfmSqsIsu8IWlEmAyWeuyF9PrDJOPh6wNlnNJKiMoFJobxe7PcKC2zc3F
AfepH+xfHwtp//1IviG9k6NXFCE6I3kuToehFpEFfBmuYBIgZ4rWcVUif6wimhGqkryP4NuO2HqD
F+chqE3mN5689GOWj26UIn/fxMASWmnihGMKNXqgZRhTX5X4R2K9gHKGoqUiHOhXEks73zbB4d4m
cQpORmWRk8urAQOfY6HxleREYCytTSeCaico7d9QK/HnOD8SszgQfgc7LfbxoyPH7IZVwaS2QVbr
t83cvGNjb9AH9+DT9C8nlfwbG53iglPp/Z0FznWJeFFcBZWP/ZSVQxFx093rTKabOdcDCZa+0If3
QG7KSzbFXV0EO19Pkp1p23eEl/eHSMgh8g3SLHURi98PSbJBBFIqF/R4vWCh0YG16FAZ0q5ukDfD
2c18pKGj1sFnNelSRrCUdZdpnuwkYQ4uTjtpy250GXibtQNXE0ELaDUenmBwbxZh5ie/LrcWQNIt
BL1mvVReN9dqH0WYMvIAHFHnNKDErPbrTDB3b05qa9AFsksE2/AdI5O3UzBY2J/Tvpn8fIzHIPKS
sGEyOt13YD6ms+HIBrnGIWnco+4M7LavobFZXHkdX66tVvkR65jU2oIdn1xDVqhvx5EzL8+8JT7J
xrLwlZyli2X5D0ezZKOpFNxTCNFL5Bxg5VKPktChR8RbnGLxmHnF+I7JqF+6zh7O+tdj3YKSW9Og
VGJrIciNIfsac0cBRe+GdcKyxkY11wxYL6zWzOG20yO66TxYl7ZD7+CfRZf7G9GrC9mLG8RzeDUI
wlSZLb3d0UHjl37kVA2Os7TB6NjgImtJew6sQ9BNOUX4huyN3fxA0VIIT7hC1RAlRm3LfAJHAvwj
lvoraUBKro6OZk0NyMr+WJC3QsT+mJlbH8gehwNCmkFD296VWubdo+Dy5S14QiFenubadVS5QoPF
0dqQ70mmy2g93dtFJqGv07yLDrY9pWqdoNXiXD5RdYRUrpyNt39nbNDeHFupuLjOOKOJpsywuBcd
O6Inr45QtFdS11XeDh8fKE/bMtjnSuex9CrNsIqrWBVNZ1QryIvDUDOGD/+oAOOSUkjuUJU7uj4d
s5EANqEEaBRt++ZAPZ97R1V+V0+YVPSr8K4v5lJOGyzsocyp5znr7ATEe63412/pEPjOmcf8YJWR
dPuZ/xBV66aU8NGyhNODk07BcowAA3vGsd9DqfWf+cBZ2tJ2rcijFMuayk9xEHKQe3f/Kk+p4Z2v
xDIrXzwtETfNZnHnIpjrQk7jQP6hPGSLea+8eO/DV2WzHe/nhmtnJDhUw/3HaiRDn3eType/f59I
1fVvbgBIHKrkU4LU/9qIwzaurlmvoUOGG5y+WeLtxUF6pCT+IiK4oWLeaox9zzthDNM1NFRdh4wq
lWW8GGK8g/0bD0aKh7aQ9sCY4iDcVKUyF82U2Tk3pr/DZedwdiZJtlluJrZEHt5SWWuIQm30Ki72
GWXyosyvalX5QardC/wjK20CB29EhszMoTnSv489EDUqscAETPbA4eHs4w3geaI7kfLc9VuKvs34
BNpQXpA7ozWYS6LdOCLtIhsUlBPjYzedIR1YMV6Z52BDoaC4ZdcSxFgYVRPg6q/81wyIaB/4GYqu
UjNTgAhgodk6LtWcXNdAHX4CIjC2LeuCJpHGyq8KRAqCziUa/9Jqfa2wf7IlvTI3wi3VgWJ3ZTpS
rN30acRImgdqScCorz5X0pa174/O4AMmTBftYCCDBQ1rmPtb6SOmBzg2J0B4t01KhpF+TWgbuYrY
RDI1zqdz1eNvhi0U6imIiUeCCeKIth96KNACeNyziPz8esV1CzBzX4/SudUxR7/MfBv/NKuHvQL7
70p5J/dhLK1oNx6K6uvBvqbvTp+/+TvEagCa57oIuQ8UgkoFi+nMWP9q928Xnrizz3ZWRd/2MNnj
/b0dVT85ZgqsKPzFrAYBJcA38joFRXXqMrDQX0g1fPqVLuUPyVQmWXONlsK169B2eo8mz6FpLbvq
YBmmdKzzg8qK/bRUqRrDVD8j0Ep1pG1KrT4rqbt6Ud2jAVbVxNvjat0fUGq7rpX4CyRRH/ZPWQR4
d+Dbq9FIgH6iIxjYdnwqvcrnfYnMfU+0N8ad9/6eexDlL4PQBD7VV9f9Wn9PWRq8d0LFfgNlmcAu
7N6FZ8E/orFCeXvHqh4qm6RH81+2V2LMK+SINlSwZ0WU3NOdAutK5nNl52sb/6rxDXx2VQ7MDing
Syx2a88H2mJO1795h+Bd0bhePYIw20oDxaduE+uBjiUxBk4Olx+yDVCVc668Juvw//Nyzred0S3K
Lgn1tqQ/4uNFiAPL3DI0AMVNB1SHPlAjq7dTkOzmOGRNxpIPut6AgGOPgN50EynujGzCP/S7gHm2
tp5/Vf5rhA2G2OwWAJYNuevnZ03/aKLvXfitoUPlBNxrWXdCtinrwbvs3LGA+i/XuJ2u6u6WwEuM
l7UQl7oVv4Gag+MTg+ZPM5ybn9iEDGmrjtWl0dupOKfTL4YkgCFvFuBnT5U+1EW528/Lyz6J4Vek
wWpFju8EoiNm1G39fhLpF6Lj8A2Ur/rsnOtkYsxA4dMIQg1DfrqxH//Lhzuu2/+MbcFjOBGG/ngT
q3WhLRI0lzZKv0oR4SHi3eZ9ufpqwCvz8RE2jxabqxHA6GRS4VYT9DToLduxK5YUNce8nnBfNEGf
gJFoPvtZOHgDVHQHyMXtWiabiXEK7AfKb7E4A+JJA2J+RCpCZwEpnLm7rMDUV7ZRd+HXXBxpIm7+
13oWUIivTtuMvgMLo8NLw9pgS9hGxibuu5/YuaGsUmpWuwDif5l8jzSkfXTXkIBnpetWC0Wyn5SG
Wt/i3aF8N4oGpkj/Eo1Lonk9JTvlaFZjSKkKHCre1rOIwj4MS2e/OdWlhQAHdHxbTdiRFDqE3mI5
1WbDEvIvkwA/VUtn8TqcwF7N6oN3cN2Ds6nWJVXK1VUd5FLXwPj8N1Hew+Osv3tp4AkhH8QCNqcF
V5Ki0OcGpcEJqEzLHlKrZlNYQPJ0ScfaSFk5CVXv7VmxnrCkQB0Vm44YdVJNfdAMULQSW1fRNjlN
KfNRLk7VCXCYCs5JyOtLgW8/8FlC7pjvU0rN0NrbhLE8aNc30/ogzZHags5+8BdyTAW07W1Fvjwk
5kLdmv7Uav/viS0Bevh4AR2lmsJatk809oo19LtwQ13SYsTJzH/87JRELCGltDLI8L1X8pcyYDMs
uH8QszbHJXK8BAcIwY5JlDhwORV+HrKunnPXmxsCdWQ1+tEYFwDm8s5UCFtFzfA4RfImxfm+uB0N
mVHCq34RpV7KbDPl+MctE+HWfye4MAwi/bNdECqUxIYTYXIymg6VQW31+xKQUhOgBpbOBQX0oCGN
d1Zz3zgMsstYjwVHhDboqEMbdY2z2LZKYxRknttEbUpjv8kkK2kZGF1usldCVW/nOkG+44/Ps0DI
7plul0pqMqH6QS7Z2eVG88h6ZdKNIeSZV/1UqBf4Krr5wGBdmbjQ93hqumB9SmneW3VxScO0t3jG
4S3ZaglLw0Ln5uB56lfmhhOjbswNt55MpxxQNjrXMoPi+8pTHNZm0nI71MuhnCXd42uT9l0va2vq
5TeaeSab7+sZ+Q7pp6hleE5jRmqlf9VkSmiflS9msIO+Mn+CdQJh78Bscq2XG0CxSpwHJhs0ZQJD
na2+UsIJg647iq1VR5nEQHPpnT9mZHGdcFOG+VzJfXwPSvDRpmWom8QEph5gFfoKX856lgHbo2ML
aIegqDG4W82Vn+HDqYEywnI8G3IraRAU3g8PDdZjE4Nx8AFZmwGCTo3SMbB1pevRsSHLUU2SVQcI
EdRg0Vy89+DqUNAfd/Zo/U/78/fKCD6XDdEt1ZBFJSvNrnCetzjzbsv1/TvlbOAr4Zq3TqcPwC+n
S3HI2jvas/6D598QhAVX6eLeyg3jQFnZqEpsh+gTKtMzIyetgJhXpkBZuj9JKRO8UMBVC7/cJ3+I
9eG7JWNX6IUymY1F/cMz2GD1A4TA3p3htZXvbBee8hbi407O4k03rz29aFQjO6BZ89x5Z0B5AA+j
iM2Ap0Kkt94LmuxCh3n4Ip/KJYfCz2Opd7bZVKQYKp8ueRoU+XNU8lmUoIEeRnaU30zOgIYIsMAd
PCqOrzFnuq/qg+6di9PjE3AdpAsCn8aZJ0nxUYp+unPZtX1U2nftFWm3mliw4HRlQsWcI4GqOBE9
UNqy7VV19qUQgbB/HWlQ5pUJm4ygIX4JJiumhFO64AuNvRvB5NDDmqCf680QDqwbVLB7PZTsfQM1
FRpoA5alExKiq85uL/WYImQKb8M5WpbinvUH3tZjuzou3D30IBobupG3JMbT9Zz9WpbZ4YFeSC8t
yVVu8LYPOs7bhjyNGqCdMxqcXSOVhDZ/p7g5ap68j/XDlRyKTTIzy4banmw+7eBto5BYYc1Ud50f
9RdX+VSq5xCjX7VlH+n8F/8UNUhfPHoG8iLNoiwLl3+mbAN3BjEnQr9NuCLtKe9Y1q2Vu0LTZJdv
5nFsLRS9GGBtXQbbakYvFxRN3uAPKhlO2WMhZMTflLRLaFPHckEKpY9a5d2Q8H8BBV+jQJyn5RxK
r+W/MGM5YOTUn0VMqQvMLMdLkP/0jy1ndyq94B3rBCGcXeb343yzwgcbG2727fi+4GAcgIjP9GNC
1MclVHZIQRvsWNpnrzbBpS5zO2SGp46m7Ay2qeWNSgYxCv1noVGbrNRoq3LpjAmhR/4IPwhfYwJU
lTuPZSZl9kI1nPfnz7pHr2+8RGfDjLxqf0PqBoKZV/QzAvzPW5SsIF4nZ0wBjuO5iWNT+kPCj+HW
dM5i7DNmRvegbRigsj8xvGzuCgnLM7wIWuNVgGMsyOzKYtciRd/R6R5pVjCLQps9o7eEjqr09qWW
J1q3ZDgrxZ+nGMwcHQOq6v1nTDcOhEbldjPvPPfUHmNyHrTetMc//L+vikH1bUOl1TrboaOt7+bs
fzbWlx6Xkt6uXppQaGCFHayKlMQ0H564YhNZ5CYQTaNCs1K9UG7TSLWeahfO6ootZ73LgdywoM60
QdKeOE1wvwm7/sjg+7tvoaTdcpwZk0YhY/tvPQd4/u9EnfjqUzdMuofFG6V/EQ0bAxD2iWd2iYO4
QGXb3bG8hohvAtdu0ECeXW7VrJsGw30OJNVkVmdeDKdr+OxZ4j2lMdEUp+WTg6lr6qmpgRXYEKkj
QiM/bupt0SfWY7dd7N2ILDTEAk4sItq6KY2uGoyV+9HcwmU0k6scbJpXeXEGT3qVGTD1mxWoX924
plZ1QM8BK4NomtD8sSUIRTKMjxNEqJHoqLvUUzixma03IfB4BDqFmnJyZjVrGA5ZsryshBHkalsx
/o5s+RIwgoiZagPh7hxk/RwP1eUdwQGP378sAsjnck9Lr/JejgGrM36KyKNSMrqRFDnlKTzpt7Yu
QR57PQ/GCuQwyTVSwaUzKWIufabKc+bRMQdWhYPnWtVQpvIjThGCYdmMNG5xRwPAePeZqOWW/hrX
7wxlUFnzNMpWqWdDWqjWra+KoC2lfyn5ozKC1GHtgOi4ewGD0f37V0hlX7e5Yjz6yyr2/Y8AhssX
9FPlwkaV156hSBzrylwwbgblTuabC4Tko403WK0rf9D8K7TDxPCSpTb3osVo4S12tcfn/mDkR5bZ
YwuY3QlgKyQuuDWbcj5sZs/d37tkjVw3T8mAPjP+OYcdkwUu6X45ceUUPr3JQ8B3OI67O5Piy7iW
3s84suQYpTjn4qu6Zax5MfvGyfha4wq0ZfKPohaUW9Qhmlsc36w3bqca8r67pZfxhrLtnk1AdYfQ
S6dPP8dVP2NPaMcho7R9M9+5wrv+1z8f+1JNdF1+xN5836hKDvOM/ry6KqgPpe/jQRkWSAroPDSr
jMqwD7O8MLaN4Y0PI+NnpBj9QmNU2vns1mteLTJ0kjiMLeCSw86jO+2AYerARSJaTyiApI3Dim8j
vI0Fau/ISn+xhnlVwShTvS0YPSPu0ogYVOiGRXqG6OxDXPVF4slJbI/SG/yk0yxyC3NK88OvDSVw
PkIFsdewTeGLmz45VmvXqA8Ea44/2NqDTJbTHQtavRUMcNdgAhxZtrMVF1XdixaeYY4xSfzlwGw5
62eq6K6CM6rC0zCi/vpDQmyxFhrJqab40VxjQU04mbzJx6l0FVYfkklC7YE+Erqmxaj5QuJ5zsaw
jEcO/jurxIzFHlgrKuXWVj/h9B5LzWOx6yGElMOZKxyHLLEOBqZhzfgZojYgcnHd75LgtBwTgoCw
dWT1tIL8yU66iFwnkvehg/FPPXBh32BumNX0PVRvyY474dPw2t0aELk5nTSROCT3BMDzzMNNUsJY
M+y3OP9uXRT7lbvvC8INig9w94de/cVLExg7fVuh5n5QhJTW740RfBCay2Oql2SfxUwCU0OJu9TG
NmMjNYt4dRJ8fRW651Y8X4sFoD1337siuyQ+0wCUACxrBx/YthEFxYUYuUIwR7Tp0Sjpmc6yLwqj
5KPc3P9y1TXMO/L7A9WNbzmh3AITcIgiycBD1JVlgwIX6v+2iOTLOto90x5QiSj5GYbiDCzLW74K
IrQ8DcRh2Izs3Q1W9x7yYLpWXFB/j7Q1AZKJtZbxqhoLQeTcYTyrl2fIdKOBsgoSAfuCYQjbnHyp
ucK7voJ/0DkcCImxG/GRK1h0maZcsEMEt1zUeqJwJcti/XRwyxXJkjqkPJfnFwDluGPs04ARRkVs
9QQIhj3jQUrxtOz7YLDZWCMcw0Hhi+PggT0veU7eKq8onJQibDhNyCLYFksSR6Pl+GOdASRcibAc
a1vzO79SAMg4Ffx5NNL6wIoODYz0mFh1V0oqRprHZ/HTqWr/SLz8NBdQjX3XVNQrQVeLX8dE/BNM
kBr2nmBIaV37GR/b2OqtKGmQO8wIK7iLWyrqIp8OI4QJ8O1JilxoFzTxI9h08hs1raQmQ1aj1sL/
D0SetgHJjHIZLdpZJLxAfIvsZyhfLI4cWN3Y9YgVtDkAdVnZ3fWzag8Ipngx1/sqexd3R3/oiKiw
Q5mf301ake2OFp2KruuDgbZAL6A+zhrgnNOsD9CQ244oOxmhyA9jXoxgEnAAtUoSWsKjVQAxIw4G
+gmj83ERF3oYSwa3zxXcMnBb3cBE501LP9bWITE3STobljYSA9IeYjTOFodnzs9IOaS0c7T2Vj2Y
3vMCncjlGBwlycY0NRB9IuX7lrVTVMnC/QdjxsNagdHFjGewUgoitAd+Byy6VjKfu1zFJwpCNJxN
pmYRVwfR4E+IAR10UPFQj4k/rlr4Rdwvz4yScfPFhk8e2BIfkBJP3Z7dmfy7iBJB4eHKq9kq8iPw
YyLiQKRIfWL1b4MmBPFSUZk2zCXMVeM2uYPrr/IStsCnzU3NWn6TlqP7CcMINffBHlGiKqRg4mEd
gBqB5JncdnBGmdGfN7Ft8+51icXntFg93sloKLLLCkJ9j5DvQ4IanJxqqx+xKs73D1ITWSc4nB/l
yxIirBpPcDwiH1Um9e+yv5bFJWTL8JGk/scKIZ7cZKwaH5uaEjg84DIXvU8/8vUhIeaBnTi0a8hj
ZQMLnzOBIDf9LEpgeTksJu2xdJz8m9gC9a0V2eIFBH4L3TbyYsGb+51VbcjIr96rBfbH5ao52YVy
XLlEL9HGb5D26FP1sN915W/GyVRVEP3qQIjPc+4yz+9exziQ2zkFVQ13MPDaRsvC8y6D8k1wxhhl
iTjPmrCsYDE3xfHtklITR5U3NxhmIFPf7KTAIkotErpLrWyCHIV6x+f7GeVM6TbgRV9EZSAI0zfj
r+qRWP7MEryfywiPOt1qeNUrJP6XcwaW0bVpR8yzq6MMAxjNWryvZTSOeMXYX/Zc6RVUcAPDWhha
nTBfzci5sXWAsSozCSkytLFQae2f6TAYMk5IDS9XzwkTy5CM7PlSexSzA0vK0mw6g5ein5DKLdtk
5fWxSSDQkmiuoQ8p4Au61Aeeg3D08Lku+IMyguk6JnyNAxhfBq0eWmr8IRr7E2a47PZBVlXoqin0
dxnjKDxK69FKgZ8aq6pYtwZnGT9PssGQiXkaUbTwVbVjZLelAed2QYNlKcr2R4kV0FHXxSyrKOvP
+Bf8e0W6I0N/RqCW41jKx/Jug7QI0EjbwE1Pz5CDjK4btOcXE8weMKsbLw6i4Ps+EbZZ6qxiWTsH
aLs5e5DE06Wh0skewjC2jfpPCn1G9xfcszFnmlyzfUW2HhaxRDsMFdhXkyFuJLrijLeIf8sfKlY2
ptl3C1Bpj5wjAKL17WJo8ecOcUh2o2893dO0bVe2khJU9NX4G4oWZug1fMtKyUMygxvjbEKFLDFR
BjP41dT/DQAjTEGFDW0kt+0tMZykS12is3F7A7+Shb6ZoiwFxwsUBq0O0cZQ9DKYc+B+uTHyDN/I
e9sOG0KkrGD2voSOU3u52RmCEKOiQlh9nHQj4Y+JsHQX1KWnHqPhsxYu3jUxHG0zcoDCpFEs95dF
iLh0ujedoLX5X5C8GX4qRxamN11j8M5+6KDqfBoWKJq03c1O2hmW6TD8lzhbtHTqa9kBW7xuvUZj
VTJDWt4CbLdg2KxoO96tVxhsGLQOFpDl5aZOVoKYT3hhVH5CacG8vLhbluh6OR2wefuzSdPAlOnw
KjsuGr8Qq8iMC2EP8S3i4qOlWzOHiLCs9DdTml1YPHxcStdK6Zn+uaQNtZNEuGmIoX9ec6J9Ih6e
r24wSnuWNxHuMqbXlxhR+tApvUnzOpZ541TzT39ELJgw5UmSFr0CzXmSBbaAroiP8TIwYXkFia/Q
AaDcjFpvzNbg0E0bfKnX0NxlAKN1a/18CGkwz1VWDVl2DYETjKCIEnqPvy2hy5GGxIfwPOc9PbWE
rBMY37PaU2a03xZ4ty/0zUmm5bAP1qQGsjRXYCrT/+wOn3OUXmLLmSSk+wB+77POZJvnFBLk1SRn
I9DbE7A4+yRSCUYEArZwdT/EsWyJquUDcG/amdhhWARyv5m7sz4cUuH96TBCb8H70nlRtgP5gBFD
WYicCWRokwez66os3x5peWCfmv73ob4UbUAPN8+sC+f7TEyBl6ixjAa11W1Xj1v2LbCWSOqlSMFs
/5KtwH4NwTmpMSbSqujc0QXekYmjVww+vMj55lvRqudpj6RjPyUPN63zd4Ut+umoEacsZLffJqJ6
e6fXwoSJCdc6Q614r9sciCcCkfxlX4Ys8E6spSL35tFk4zkTg2FtDXjjvZI3WcSu3ljiWhsYKcPg
tjd5Yc2ZA6pHRJHJjmDQ8i8qTjgwex5jVfBr246XH354PMvec4nY2coKQISbGyyA4NcrJa0fSIWD
7QeArsw1Qb3pEbABuZKQ4DVG1kgTx2NAkLj2lLKiNZ3Ce6/TAFgYIS4vTSx5CwsVAK69PGjzTsLQ
7x/jOXovPGfchCw9ZMXJVQ+QV0pXvDB2hTIhRgmf8cM//mAqHjMBz6fShziRAJVdRDvDvrMjMuvz
ttFqowIRy8yTR6RR1wmt5CqCdz7di5dQY/M6I9L1Pwpx+XX0dLM774pQhzqnGs3UDHB8Z3jhLPwX
Y2uYm3onodOXwEfQw6ORLp6UplVqR8275vP2hLOtUngNoJSWEuerCym1ABcqRBk4aoEnOj51tizI
Vyf60nY+1Y6M9DL65BCgRdPck0bzUW2/cTx5wS1i+qagUT0+xP8Wvc19262ceEWabVLBU45xL7n2
40ueYNWuyhbBhkTK8VlMUr5J6zTvEeJ4dmBsHgRc+tVJcnWCQWF0idIOjS6XeS2xS0lk72FciVII
texi2c3vrotuugRySEiFTgD4iVpaOnR3+VB7P7HZodr3pN9ASyy4ysTxFHhipvQpkUH2EtcPmneB
EMV29tJ8k71C6zeq/XaCR2QQqhqxv3UoJxhv1tNFIDWpzh+KOgFbyhpSPLhfgOm4KoUDn14SlHE6
5ZkQvQ45R3cHhD9txDEUTNf/vMfC2XF0m69iDfpCk0P/AwjxbT1lMLdBw+n8V+qu25q/2Fa6PvF9
fXijubw2X/1nmmlRwcqnw0plvo6JUWBScghH4oatVjcbbnggd3S/5JBy7ws0Bn+7LrQZPxXyGplZ
jWbSmJmEuMB34mSGNr9hSmkSpn6K7OOjE8I+LLY1bZQtM0tcfXQOsAlqA/j0N7HiCsV5Tm2R7JbB
MAQ9gp0lP9JZnsuHDQMMKINLoIiyhOAGMSxUZ0++NBjBCbcj6BabbUlNLE1y83Z+tOvqVPOtX+8c
Nvz4UG3/MK31Bvqz6PcBd4ZrtJFPktnWGG2PJtUqGs6lXyNOq1iKXxs3xOXcqeKNBGqfhidGzbB6
Fny72m569XBPrFmXSOz5n0Cbdq8MU8786WEH7tcACQRNkvu0ZvLKV1bwzSgB2VlbIzcvFcTeCIBL
grQTEdWzCDA68Aa5bNEncJQbKpGjRJrARDg/C0B9iu6x6daeJZ+LzD+4/xu/EY9DQQ1C85wEIpsJ
sEiEFOAUhcFB1NHxczkJavjRu7kzVVjlHiVP9bYabXoa7BfGJlpkJw+BwhUAkD4ES6tUazcYYvUs
Hn7cCJcfAG+b126aJLuowEhGDGFu0XjucXvGq9uqZaDh5TVAXoNENdFk7hXvHfB1ieChN1rCHt2J
sbKmDRn7TLSQwlE8t6n7yz6RXogbEKS9K3OOz0PlMH3gJwDl6tAZgl6JFBO3vOTxatxSDCmboc9y
3LRIQ/p6+JqImTdXJHRACQQf+WMluVXfE5xdH7UuT2AAG/Rr27EE2rW7mSOc3GNNUpO1ko1W1t8c
S5WN8vQBw/bZVoYOZKwOeYaU7e0Xtem0AREBa7jUjTivVtkfwyOcp7e6tY50N1+y+IAtpyb25lWa
5UsK/YDSHfkMVEUzLekWKxHDa1paVeltbI8w/XDxbcWUm8pr8gG8JES3H4YUGNFBZt2ZApo6FtzM
OTRltHX4Ni9U+2wj3AluAcw/3NE9Y//kvvfg4dDrsaNW7erjsrZdKPjzSJjNBt1/0Czx6s9HHQ6F
L+2xW5wo7Mx6e0NjnzIegIGZM4wWBTr0J5GOSRhVFqXRuUuZgQjDl0XGPMRSsKnrPDa7WkFZ/W7z
/Mb6sI65Bxiopd1wuMj8bA6Flv/KNofXWDe04z/8VFeNYqjXLAY6hoRc7cwICyVVOWT7i8q+CfBk
lmJEqZoNvb3ekAk8F1jyil8+6/fTPjBEKQQNothUaOxIBqWVAD1krF/ctzbbv0qUFLGBkaVFE0Ze
62Lr7AYXh1peAamwJFfmmEyfuLbT6lDrJtPhIrgGKUHGfKJCMS3OqyE2JhBhHDlMH3RoC/svTJiL
ofLcweMj3X4UoKiCWeFfq7U+iV4pVwUt3GawQ+uP80a0qhiWTrPnVTrlCksoGleNuxG7bvyDwVX9
uQzFO1gtaFkhAUcAfgC7ZsQKfIKIkL0LffgDYd4Bdl7pA224LSDkYww/1d7Pjs8UZClqza60Rdb0
ysX6/m8eNTg/6oMP5voVA7joVYVq5kYabHU71tiMnpxbKga/WqnbvquIqXOLJUGzka6QHTcEKT0F
0c2WK1Gs2hpLflpNeUflu/modUmnn7XZgyV1cOx8KZGHRnp+EZ/SEGY6TYe7zaM8F5UO2ffaWk10
fdjcy7nObgGxIvVU553aPIp3Ro6Zme2rn32x24Hr7plv2VW7CqxM2VkbLJH4ZrcYT+yT/U3YyxP7
YvIsQP52wBErs+YA2gFIV8kbjcUhuGbksdN/pxCV63wGjM09yqxwv4nHeieFqEYyVjpZY6GxuH8Z
baWSm93rooOxQbnCP0JDSjP2BIke19I5OmkhfNTi3uE5iNSFkWYRzEJm79E1GItvamAhWGN8n93N
OcrqcbJn1fXzH7mLN7DVFhRHzOl+FnmX+DnZJA4oTR7RcKpc15SeEB2FktTMX+Sydjy4m8kGUf/w
sIiQi3dS3V5dwrECDCoVYNB327An7UQ8YOnq4TiNgHeBzzGzioGZ6K8W1aZEUvioJVevZyU6ez2O
tqGkFBNLd0IXnv6nKQ9QaHIElKwTZiDb/rPzklbUnvQigSZfBd1K1TsI1jmJrFnIXhu6FqsRqU0G
sDIAe8PT7UePtzd33ARR4d/NbZns6Ygcmok6K1zhoB/3pZap5tMPoTKoafL2IDo2vNpoSWIvZh0j
kyEN8uv7rTI+sXyTL+DsDa4RSTdz3/JPBAr1cODp4C9m8LxznCDW5pn3uE4KaECB6nxaEVyy4Ipl
/T5lhnFfbzhwJ/XD/ex8WLLNvRwjHTW6lTQfDCX9NeUV5cf0LktxajZw9F1aImh3827lKfBJQqrd
GrWxotBWNyFdRO6t3stcOO8Lov32zIhd9woiMd+EvdPW2DdzC0CHjr1FNjNGSi7dewxy2Ny9nzdn
f5ZVhD6tOcjIbSe2hYIrkrkzJeMC+DNhMHFiD7C8f8cymuVsNfmfhYnwSe5XBvOKLRRzLrEFwjpA
b0K8REpfUw3gphGl35cEHxBHPj3toLAXb76F6eey76miiUDH9sH+Crk6R4C9BNhA9eqj6ItCJ503
XxrB9mzGVh6z1MXToN6/yR9Xb0XIKOVymLPbtXfRfduOuplEXVToBvK9bKbKm6FCpn/kqNNw3VTK
VjiJWJKrWOZkz0TfreTCbztzrXe6L4v6HY99AGNat/72bzQnnvXHpKRBfM6n4qTQ402Uvi2/MvqT
dG0v/SAH1r+72bzg55XHSyl/DRbWegprZSsdQerFxxdzpDwNn4DnPvDBpX2tGpAj/0QGwHFvnAAN
2cwsBqL4+4e5bJpXn+w/QnCDPFNwdI2sCAuyXo1XOnFIDa9FxCX8tT2/MexULh8XPUnjG+XcR+JQ
uXt+G9uhwS/6d6B2tcKgBD7M1rM8X+fHK3Fg468DL14RjwXJu+62WnTGHphS9ijao5duBvH93yGJ
Pe5uiUJ4MVoA37ZcArEYyGso3TKvWQNGRSjCxTikcOL/7D1GDMF0F8PZUuZ5LBQDDkUsg7wqZRAb
gFYv4awM4sFbrMtrosEg2fXNt4sUGsM6s9DshXcIW7HnzLsAW+xeAKroLrjiwFyAPPk+LUd4L94m
P2U4FTt+Xgf1C+DSVLmut9AbxOxBG4dTyWao/znN9m1oO9aLvsa2msA4ZPM1g2DiaxokvEPuXAiC
FJSQXNEbFFeTZTX4CRCPxa+yByMHdhJ6blMgjsuB7V6ejCp9Ken+N8GYMblQxRpoJnFwBVDlx00i
7o6jMzCoB/xVdDzy48ysasrsBplDubo5HAlTk1mEBq/AMKF6PZSxNLaaCY8/8MoHoMksHitRN4DF
+JGsdvcfaEeZ33m/Q97YohV8+cZnvzrQCc8sook9x9/ALUIaMYZjFWBCoWUG3QmNQ3hRU9a2RJ9Y
+N3Cp4oL+GtQ0FDr6H2qMRNJKU0Wa6aC7KtLMqZyHrBItjsC/RbA2VNJmnAnnrxJOMO/p/2axZcL
MeoihpM4p5eCOTkjBKYina71//HuRyzzt+Cc+7K8AHIiPyf6Yu0UteGTa0MxsvY3L3ryCjlOlCFb
oyQH6lfAr52CgSqep1KX6zHMnIUPdrDGJcVCKSHXJYKrnytVmD0C9ahyy7BBIH87P+5Ngb20VqCU
6AUjSyUH2SKiGDRZnmXEkh55m8Llfa9Q2AdJUYVI4vzwq9DavTiugifx7CBba9xOWWgbPI2TN5or
vpWjG/K3yddpCTYxO40P4Llz+PkvFR+GXKV900O2LXGM6RFAfJ2EqfZupQCrCxXsB5Tmhpl7NLNs
7ATvmkuyy16LqHau89QEJI2gHKnE8MGfJMzk6CMXBYZXl3dBOzEPL7QnUa+z9IglWxXVzphdjBS8
dHx2Rpc5oOUP8nGmQTp3YePm7xARvCtXhXx8+qAMwlStkiIMi0QT+0FUmgN7mwNU4AqRmk4TmtWe
MJind8keyRNoS3LHd8emRZP7rhO8K+/kYEVQCQboa/lha164JDnWxs69bBACASrUbIqrv6L/DFiC
8/tFWfPHJJOGbxEwYsVyoGNDsxBOl54WBZVwGyZw+DFASR4YjE1vLIn/bJTuSf3E+rrkGnd7ATml
a6eqGa9JCSxz+64RPiOXy6xjtqRV980ituB7fBf/ERjtaI/FAljDKXG/mqvZK2BciIXMoTdUOY2U
xnrRL+TrVB41CIAQFt3XroOUN9iTopTFuwx8xH9ExkN8QIzK8sYimi2Cyy3Mda8r2w+eD3s0TI34
hPBTqTssqR+5dIjW1ASA98fqUIIb+2zSDjmCAcsoIFCfzm8d+XEklRFb/AMA3Gi35sf4wsZoUl+1
5hliPBa81w3GOuo8JKmH5FldRqVU/vSjvaSlmwuvhh2bMrLlALDQ5TTSvUTsKaART7vNAb2oVl4k
V+phZ/JCh5gscDorCDlxqgAmDSIvrG/YNzqZk+o8AL4RZ70kf/3j32TfVcGi74q6Jeryod04JAiJ
ArJftPxdbsSgQ/UZqvLJAf+sr4t+0mZ4qh+lgzca3DvmBFZlZyQQlkEeNwJ1RKJR1BWuU2PjclZ8
yxMUvPneMsnFiQTNXdjq1aLy15sI/HAr4V4n+fZrXeDD9LFhze1F0VCrS93grqPFeEO5PTG7z4K3
4BUg90uZl20MUfWUR+raU05KnR6of4TQigmrvZXfLoiFmQZ/G0Y/yW7Hc2UR6dI56p31wKhyyD5m
UF3oxo2zlaeM++3aDTYqtvSQnqb4drFkN4P6k19agtq1TOAph4Di47DQ875kjesp8E5EoVy3ueeO
IzggFX7DFaOl3/qmqAq9PqNJRTbqq6pBy4EQW1LVZgnMf641zktsWIYsre3ipEEOX30qhrFvQgMy
plgDxsNpEqhKka1PaS82meG9iLtaugCcq3R108j4T5SMEDC58jop+Ll0l22ed1xaWpyadd8vERy4
beYOf9hnAjy0z2s4i5SxmmO812Yu2t8ux9PaEDOs+lvf/ComBt7N72p9BDYJ0lMQ3tQs27ZegfnI
s5cP/mIkQlQGupMwzHuU6i2kceqJYM4RQgA+/2sBwrCcaWgvBrq4MX6NGAEl5Cmx/rsCzGiGWM3R
6gB5q55dfX0eHKeAXjcA2hV5KW7DFo7kWgAPaCh2tL1jgxtJnzbGbPEI8b9n6SJpIWdDWr+jSmkq
I98552cNHTHMe8ZumAnlr2gGjDNJnisSJTZROVbX9iyV6BvekGNTsCPUijzD2hZISUWq6PJ8/Ru9
aTQh+SmP/7B6HTFQ6FEmxrDxujAyNku4OR88EIXOvsuUQk6T5N40ZgOH6zrygWuqcXIL3+F4WtHN
0FDpbTP1S5H1voWplC5vL23hxkORrNBhnQe+2C6+yhdSLZ4LrH9oMJQ4fPj/24DNNfqvon5+qNDT
TpdTX5mpfCGcCaZMLhIa6Cy6iMNlZXDHWOqRvg9ncRaOf93qfwRdAA6oEP1jJK67kzYe5DYYGMxq
GSXK1UGSIq9BxmAfWD1LVFyCsdPxyUUlVgQQpIAvlcC6iV/mDBXEhfjwcasJQg2uNhXFbzPed+eH
IHlAlXse6YBsV+ERuU840zDY3wcFnNfpwI5i+yKBu5p2JeGoUiNxemXyDNlVGagFQWAKeiJVTdNl
NQRVZXNNtIH0+C4o4WSxH/cf4e9oa2hhT5uUcLDxD9dJkS3EEBBhd4q3kN6OI5g7qflyzjZgJ8ri
a4Geut3XJyZF+xcIu1KM1uyaQ+4mvXauvl+Ac+wDkOYt/0QP+BLOocOmnb2kbZJcax496g11TDj2
lSgGej0VFCZVGcc3S6y9AcE7XePXeb5F8XKl2nzwQirIPcajbFng1R+Q/OaIG8ZUMDeXOK73jgBs
sxCZFDHGBTIi//8xvvvhSE7764P6Naucv2sWDuPBvzaiY/WnRFEpRFKmEPIdnXpkenx0IEqGY1H2
meOALbuaYwCleZOvCai0zRx99GPoAO+yGqAdSJu6wetC/BC6y7lUY5nEQ8bluIxIj91mPu6oErMR
LLlwzYXpQyHoypgRMkr8RvTvDgcZq+tfMyIiWYXyhK3753BMhWuvJhRoRgyC7Borx00ffSQbv/H9
+R/oE//SzDXBgKsD1ptuk6l7LTWoZUxvba0XBPDFF86nvqGICVkYKvfbG0ba2VsIfjjNhD+GcFVD
mr7O8NUSfCqcGaazqparsWTBGTo2YDnYOk1mtrsswVJ9gcja7lgV4kvgozdIHIexBGk4VHyaxc7a
0wyyy0T/PQuzc8GVzX3SEHu1Y7ZW4nGfBe9TTLMZ+P3YlXl8phyk/v8HFO+0vo/VryCzAe/U/gvV
acPWByteA9Z7zzy8/KziP4xzsBef5qO+DPHBesVmYfBGziSGCX/jHDdWJU8Ibxybqv+ORprORb9e
ROpSdDlvx69iBAvejgEv0325KFvnCyGIGaN67MNSg6HW3n80JVcm9eQLr5oqTAY5TCqtuS6WW0g8
w1hd3w2LetFm86864GjcKQ4I7n0OWzN+lilw0NQ69PPny2AOjIC0vVXv/5IibA5dUMays8uDyx8i
vc/05sFRnck75ON0PgkZFYI4u4upuU0PKpcN2aq5zPo/4ZZlDBwNgDmn0djFTT2TmML5OePJxi9w
ComLls1keZYPDTX9Afo9pQ7E2p5PUDJPm8kPl50i4o31aMPa7UrrQ+cZE6gH/Xb79cxr61plfjGu
CAcxFGmOB/zjYzTYU6PVwAANY9fuNateJAOP2y2AnDAPejUrxnmBQwiHqwktHhKiWsUtONE7NbDo
w5TWZMmdmcABvka6re/qsu5qI/U9pUlzcMqHn0CWe9I8cA9NHtO5xlsSfMFoUqWuGTToWpSGm4qv
xRV2KDW96G2mjwBfr5O30wgQlXWA4O3IChlBXr8BASG4WcZDnLfCxlZ0yTnefkZuRWcPN5qRVrpF
/R6XhVCpIiQi2isJd+pVcQgpGJyGtYxHtoO5vH3ZvdCYflUoTd0ZODMnPTuAeXhlh7v9zwoldUEL
27nRYksCWW/F+BdfXn5W6htgODCaBK0R46Zq5gAPVeTy9HN4YsbgQXjHmTciBgl0JyWNwnEAdKEO
gUmUh2z0m34AWWp+fMvXIXyCe8XpNhROosjirlqFyES58PFkAhQdVct0+iwWwZVdrXhpeaQ73rc4
36z84fCt4l4wU7/+WocCxrEA+5hPojdogJ0DG86zZUAf7PrHmTQQdVBmqw+KwE1xpHeRvt5qPykC
PmT05syAG5Qk0B+m7lDkDXAQkG9fvBZA0OmBhaBNKCy+DqHZf40uUCMKIGrOrmHSjpCEUqp9POW8
OLfR1a0XoaH7hC7jK1szsvJkce3VnVfINuO2b7v8Q/rUzd3Rt05ct1NhXBLKNN2+9TxkZGiWMywi
OjusA/am6MwF4jVnkedzLymch4Dum0tKRUWWRk40OJBF4n7c16tt4RJEbDT1ysILfTYp/5003BIh
KOtKSo7n9KXVEoabHALvcsS1E+69jBCBRQZnWnCZ3yBTvyj3IMHlLGK9tSHyVVZmVmy2uJnWr2b4
ppmpv7pxa9cQa3P/5cfsORnm+TQCWhHp91WHPq4h4KFOG0TiZmBJvybjlNvBK8zf4EmXfhCvgow0
NeCdisGKWlyxYyEbCpHetNUXgBcXqt+uLmR4rxQ7LmTa1VQJkLwdhQ5yU1Hd9Etc2WpNAKfLwiL9
ZsQURn3CuJQWqN62CdyMp0+07l++SWzAVxg1+dRp+MQv0hAbZnzeRqNJsnLGzh2BjOrFblxDj2m1
KR9b930Ise3J5kPwlZOLWQu4hYeR5Q/g8mwyvfUAta1+Z8keB1Ob0SRdMz+faKbGS9eaQsaIOJlT
RuyVcjb8ImLxUeuhqdW4I2nWqnc/JtX9Xtnp0Ua9CvSV/A4P/fX55ckPWqV5hJ+cXw10BxUJBnla
tiZ8M2bUzHm7EguUQrFjwrjkQOc9CHkeIvolh6557SedHa1Ckp33B9pJHNWjqHOhd/qpZryD3HUo
3E0B73aPMDbI47mH1A4mRrR0+semh0kMt+wY1h+JdpgP+gJnPBpD/yRCrZdPJBAMcM2iGSO+2Ity
eWhFlfTt+RN28XNRYZQArs7MUHgxE0o8YwXw/HaVp2/hI4dVNZwQ0vTmWvgstD1+uaiMeU136LfD
ATxv8BQg51NTi1scFy4wVh19pgI2OlMY9NuZ8euCAa0d71k+KFtDFflSOA0+2jo22G2JlUnSS+ve
C/pkNpG/d+xDeoMcUrfa+a4wMAEJs/sJ8SP3v3t6H6IdVVuJiAJ+9KoiiYONQpt/8IcQkY0qTlwp
8iI0ssIbIOJ2VFxssPlq3SrwW379iam5RoefBAxU5Q31H5LhSHHYo44UgnhZKezpPJtR9o6TmjHv
K/i5V6ODe1cYOibfgbHGi6gE1rtV5LeoGET6L60uT1nlK6Oib2GjQx4rpRWKZnqfPMfNM3G4ibHV
1N2MnAjxkZ7FBr6WKyQO9KysDkBtbG21HTAp31QUMmedi2KukPE+lXHqzNshTKHudIBcKUboRdUr
ACToxNBtz48lHpPC7lWtkdvkBECjoSkf1ykSsPkefg/Sfv4eFHXHfyWtyp2iXIAu+281cOwl4ljJ
yS0RlsKtfw8MuYKyCh+JfxTjaoljwCtXRcPomT6qMupeXqEalTry0HTSRHmF2E03lV8HinIJaMhC
edUsHteH3eaPQgEemWsQ8jNWlzAggppWtzTiNVgEPdpqt71cj0dVz+0uxiE3CjgnE7GfWZ5NaFrw
mn/ZkpokOywkxBAm4bQN5BNg2w+G8+Id2uQPC4Z+Xy9rxGdJex406LEUHmkvE4XKVWlA4UwbSAP/
uIx5p/L7vw3T9uxzTspzT7YNlpYDg6FDQYp1d6eFTe0ISRNKtyBurFTpkdrBC+/k33LlkRJxf1LC
WjLbdekpsIA8rZkJ8xUDADdKtYKZXPI8inbm7k4xts5sQIHMZLwqcDWdLPnWsRzGMAHHoHvDChYV
QOn6w7XXva1z63gnRTo3on8KjFcwzMTlKsSI8xkuAMUrsEpiI75Up3S1+qfUsKGd3b1z4f9+Q9Bl
dbiI7/9h2oRnex2/l71Lz6qiP2kHmqxNTg4QehnefEdxAQEFv8bBzWExic1EgddSob06f8GCqoKW
i9itjoPk4GDdga2kYnLwPiVGWeaYR7stMacL+9IlANNel+58kw4KJ1flURoeQ9oDa+On84EJOwts
MxM51oDM5K/Aw9Rft2pNy03CZxvEpE4vs5GRcd4QgSo9aYNM/VfDpKwugss7ZoLo/pfAbt3pbyI7
Bj4pOvCionP10PsaYEJhMreN+Ye8dir7WagSvWWBrD+MyuWOGby6fjoM0hsUahYbOLepNYB7axTV
P0rqBDBDzPrEPW+5g+1Ku8EI6OWOjEUV2bGluBMhpisFMcf+7xs+SSJ/FRjvw22NUBzxUfNh/7Y1
mXfrGCIMCWCXFIojZxaF8sgekSbN+IOiYaIqZOePPoIVZjqHlr8tTPYFceQK4hk0s7VbTbDCb5//
qZQdZuqsKGA/bnI5KS5R8KmS/AIXRL56f6Q+yke/4ZaDcJW35fonLIAHhp4onDsbb+rtCgnFEtpi
0zRvLLFJR63licIMlQo9BjRijoqp2cVO3TtaynrwiE5hObRCJ9ne9d/CONaGdROpyLlOMv4uiAZ3
Hz3098k6NLbrcOexUdpwDsPQXZftvUQwNroK29ZYPxKNeQ5YJXMA0jZgiKgM/ukhCG6YSlgCqcbF
6O34crngLypJC9DKtPpgTvf4HGH9scGUHjPRmForl6YDcaiqomuwlxbghVsJy2TFXvfYf66r4BDK
oCLjjizOW2Plnx1Q2npVeQZfJyogDfQkWPDpdJoQtQL3yfvbi2J89anYmRboOnzMh94BRvC0DBb8
DjjNKbhPVnVLh6RVsYq3tsk0aIXjBtIbh+Jo1BeR+eRaC6hIywGo2RFKl2k7sCNhCEGfYHrGuWEM
LwOLG7a1My1Sz+Sg/+7fDwFZs3wHaZI6c+1hqhHguWGZFNoNlCjYLfl6gMHfMuSuh6N2whyXLQEO
/7mCq8lxr5AdeK/0AGEJgQlxOCHdTx17tR4AcOBHATNg8Oy5o7tOL3vEr5ap94n3l0q+bqp5HGs5
6KMx5Ma4CC4i5u/ON9KPNQumuToWlQTD69yRnR/+pGpZf4jBgx+nE1Zzn7fFA0bs21vjYftfiMFH
T+HkkSC/uReamf69gZt51hDkph3C1Qb0av2Qn+C3UnRMc5ylX2LdrRVnCCzMH3RMrauHM4kNCCIL
ARI8mJ450Wakmrf5P2THyc1veExihcjzA+8vCMy+ALe1ejrBq+RXOh7ODuhZdqH1dfyhWw14ybl5
moI2Eilcw0Khjc6TrfBuyTYjdsEsrYpgYdpfptNxrwgQbbCJnfnc4fV1DvxAgenwl+qy/JjVUcOj
fKCvPy+xXxhBHnTt8+y6glCgvZr7JzfHAfRWGvY9Usvfxa8ZhO8Wn1fUXlr4xLfvhmVIXd5Lld41
Z0g1frxwz7Dr850Iyjs6NL33ALNSVkg3SQ2wdQQAJO7iDskCNB0x0HfRz6TjDS8T1i2PoRavNipn
Z1tTtO5p9PASsJQ3Z5z0K6RPbNPRR8fTML7d2KIPLE70+NngylJPFqQDoqfZBQHoWCe8PCttb7/5
z9uzTwltREG5P4Vtmx2Fi1Hv09oYtIwogwHyNs44VlyDcBl9Mz2kbXEtGjpB4DdHYgAcnldcPc82
gj6J7dEdEicekDxe9KhhHzfHM0B7QrxGHNud6BsQlbz87R98o+u2+rww4RhpQhvTWO6mCFlV84J2
7qGv1wbFuimTlWZoWHCH9zX7qOTmmrtEuNpROXnQ/9CRUoI7BgARGspCeU9/DH7joekA2kH1v5IC
FDED36aHOlX0ZCMskFpk+COMxJfPaBS2GGn4aljNvzlI1Kye4RrlDAtrAwisptjDd8oYdhnYS5iS
ty4V+HA7kDhAdGQM/VSmCgYJtAiIbo8i2Af8xldsudm73WtE57WvOKPGF4eVNtnxNcfoc1q4I34i
TTIVvv4g4hnLdyFQVO4ZQbGCEWZ7un2CKzveGa4BFjnpTjMTyPZqdqfpYGZUTetuHdMatyca7JRJ
fUdAMzLLmKdPkCDliZJvdqcUMgmNI/fksXQslZnyHu+0lPqGQSIq+aeSzNmiI1qT+9AwpNq2E25s
Jd65EBA51acub8p/Ei/QKGrys7rjHBw+1xpNH+Sjfb0jc00UX4+xdr6nhl7t8s0eVk62DjkOVaAr
ecadXRUxH/5FXEeo3+qBuRjU917XQWG7iRKqoS9xr3LJI47CRq5grtMNdx78E9id5W8Fl+JpaYFS
pu1sVOjQHPhf3p5nz648j2fso221xlDgKhu2imFwl7xCBqq9YGhoTVq2oiHfqb2x8OFl8cmSm32i
UtnrL4InSAuLQDSwHiI+Kaopjo1MAcXspmE4DYVBqNrudnEJgQy2Da9+gt5bItx+/u9tjXydDywj
N495kSzqvPPIGNWfWowVSLgZEcjdDkRCaqEZSqesNsxlvIUcr5GVPLIu5Cz+RZdhMtum+f1S87/4
YKa7nGEyNLhYtGLxkQvOAVhUvjch6d+8rPYcr7ASPFQcsGv2h7TghXlL6DcxGg0wsYG5R4ev+jB/
XZb8k6UYhv7TsBza5ijlj5mVo0VQPyhK9hLjFP6HpZnjMa0vL5KGO8BM6efLUzv5Gj5F/loOVg7v
4BHKBjVqgi+kP670RjTC2gO70YwoFmwBvlnPOdQmD9xkpwl4Kd2BHC9J2VcTpPM7ok+iLihX34GU
mR5mit1sjs3U/D1J4FDjYW3oezbw8tOciqMOn4zoXkX5wAaKxWgbFH3SKQKA2peLatlFHNdrDJIt
zl89+93eQoyhEwH3rC8I5nWOZMX0wYyaB7YF1XxrmqTLjrT+FpbNtj6I+BFjjvMexSLfMboFdN3L
jf4zQFPNLoYL+ZHl4cdW0uelXwz3aNQUAh30ei967eAsuYeNDoFC3c+5OoYtpYLgYV+GUZjc3E7x
XYrzYqTvXgdFJMwQox2AoE/ccl15wfQ/9Wr7Btt8pfb/aMOmiuZSg9ABovcc+pIzfUzoffQzR5Mk
opo57544t8F4x1SAURBrtTJKcCWs5sc120KEGInFaXG34DPVzt1oYCmcdVP45dsX+pO7O8nJ8IYh
rvkLVB4O2PZnhZkw/T1R4hWzwi8ktsgZp9Es3TzBqTAVXltv3zqUrcJ457xEOWH8rpzmD55gTLU4
MHI086d2E2rFAehoaI0wnjrAl89NJl+rstTwm9bi9TwzxTOU5n4U5iWmSsFKCY3id0DjpPyN+5FZ
4dXV0sAP2oHaHG1iZd8GxNJvseoFdnaRJcu1cabW6nnn1uJjSs/RM6c18b6zHhcb8X6T3A/v+vl2
XSmiyqIrJxp/qIvcsnPlpnyb3g2wskqA+8dvB0FdsYkUum6AtdVc1eWczG2bPhqpxcALxpOpHtUM
LJr/QKYvgsFFf+EgEmLqPmIlajDGxCltHfOsARlUKtyEjCxyqwUJheGWVbPXLi1s9IWotSpW+PRM
iGG5KjRaKYJieqxYDQ7FHc8Kg0DPv8zfcPZPZqrxqIEJyJSff+D13RBiVcW23Mt7RTNcKNXMc2xq
vt2ZUQ/6cq56r9hNIeddBJyH51O9j78iGur0HtOVTsCy3GzPOdcb/3VcfVafaWmyZVy1exu1qfvO
3ylgpwOEH1c7I5jVT7pq8NoOC7tP/ZklXczzIvIo+NmuVnrlvGoesuNcEdZkklHGJ1U//Q9/lqLX
hruD4mHLft8+D1IKwSUdDl86kHRASwaMRgThPxcT6KnWj1t6BsELvhKOongS0s5GKXKLnaPSW/j7
cpy2UTH/nrF24G+DUodXY+nZuvo1LewW08q4JlAQPHVAM2y6NCWE3H7b1JfQg7Q6x4CvZJNahEZA
2c8I7juSwJBru8sy+Zg6hxPkuvD7oRIFWx1JMzrUDrURR9gdKDKv+1ulb55dWykOl9fVSiqRaK4Z
KF2B1QX7AQzc5L0qudTRxtYGk3dheArem8fiyKaRoI3lLUN1Dv31K1HXTTfMOuS/mONPkHQka6O6
WcT7hX7q8JrrBsu0532MrJB6j+huMX1fzivykm3wI0RziqcszLWSobS+wfaGJSGg7de+vsw6QGSy
8LpTJNcXyK1YbkSCA8zka4mioMw0K+koyGjWdJYJYv52puo1l3UXyD9l7cnMJdHUV4KxP5HdUiXN
Q8MyB1t8XlVAsIxZdQgm2QkEWvbIin5DYEbm16B+b8OEB+Gv+2FHBUplWMyfIHHy4Vf1yEiqxmJ7
RonMpJc80oQFWBTjapNQJxtpw+/alivVZ1S+mKxz7u7itzyTBqeg23fM0W18nyusikFl6d51D/Gj
r8+gS5Qcft0+slIAzIWpEQTxGMDeRn3DPsmoLzr28CnLYBLgIr/fdMqSklaabhjeo5agsqLlWsIf
98V3VR6e80BSTzHFOrSkexMRxS3X8LnIxr55evzA/99S2+yRFkB9yfrg5GKUCSD5kEj7na5WlDDP
NclTokSgm0xFKdvnjPxXjIBskMKW6cULnbSZM1w23XtHMjOKWdGleL9cbODKEq7R//a/A7J8lzlC
DWOO6/rXyCWdYqFtsoAFP+qPAEvwqET3+nQC++Bjb/dmPjrItLaF3zHFHIOs8XsXKAQfhcd/RM2G
fmBhE3Huwyq9NuX461UEJZQYmK9xPfYgYnPY8pP6LEygkdhreR2ZVhKu+Ss9lRosU/hjK4vhqslA
MW1QjgxSRTQiuvPGIgXreJL12X6ihzbUXpCC0EFEpjNCqVyNUQGKfMD/vzeoBUIuinz1f5/51rMX
Qp+L3yz/NS5NEf/w7seLyTCdgWvJHP1Bad2zzhSWy8q9qUi1zCOa2umLPbvc3vpsG1E3cDtn5MCL
fveetjKMqUgxS3OPWQcqBIxttHuN/DfHBwYKwdsVG1w8qWPFlTHomOvu3lGooydJfoFB62vGiMLk
UjBjh5DDUZy3OCPNgIudCVqqKFIIDdTGwdkYNXZ2dSdfkpvT+3DsLx87GM5mbCcDMtHDaRIW9Ssm
c50DIWz/6Iq+lF+lxmNQEAwC+8lK//Aa00iQCRIUGZM7AgFXmLgHkY4eBvt5wIe1YGLH8W3iQ+KS
mgbYcdStwBo6ePZVbmkEHe5NxFXtAEmctktrJtAyWQnS75A7xGmJvO0LX6DHAlSTESpvrJg/xMu0
a40+fbqGXxlqEe442MBxZBCznhhXUnwOKddw0koGRe+Kn7jw0LCwc+gDc39aHC33rSdGCP3bXOIb
YGu2Ig7+V+I83wDhSICFf7w3cl7NWQL0iwkkL4HFqN01hdWXOpZ2838kFIX39Q/THLyzRyGNaIb8
WEFm82iysZMqERgb8ozDM58Tyx2FVW9w8TslHqSVKBgZK60WoosXb+Fq7RPZ+iqCRhI1rbp5WacT
dyGUbffXQ7HewIIwmEOdNwlLlh/ESUT9j/Pg+GJrgg+YfnmL7x/1kvLXPQuCfT/FaVRbk5alSQfo
Ade9aN43xDztuMEvBvmoIr+Z+gqj6O65e8I7D4ejg0KVHYXYn0JbjQU1EcKniSRcnD939ml0c1lg
rsHvdPyDp3au880LGFwWW3UcT1Q+fAK0/argqtOCV7cCzAPuhRSLYkhluHxxU+YeJt1oIGyHF5Ge
1C4LnSQ8+Aui+qOQL8lF4mp429xaI/vm0zmDk8z8VLsleeJyqu5oanJWBQqBtZQ5frsxN3o7iM4c
JSWthIgnrR6ovA0vB0AmDQ0FtY1BorVZUVdikBAIAbKWqejJnlRhz1WZ2UNF8JmuA89ajZFGJ9MK
WcNDLY1fD8NIVbI2wACNk1d1obAuxZ+ynPqUVulZgb4jbyqzZZNDpy6iYF9wmfOLcGR9p5hLUdMh
3LiePDR0HgMgtPyT/YvQCE74pvx0AcdNWFGlEvGfWcAaPxoXKrvm68su+y6+dLhB0kX2msxMdGiu
Kr9kr1ku5Fb98u/W0v6femfx9H9SUUnWKOS/gGO/gkwoeFL1lqEQtnFBkJEv89TKlY5PHCrs7Si0
y9KFfozFhuOHqPJ7sRR/ODEJKOoBWXqfrzRaadedPC8exJpIF/b4x8xxYfU6334i/txSfmEsd93w
ilQBj5scoL2D8gMlWi5PboRWX9DJ2McTEyqxz99apNc88YHcXZdpfV3PwN/GTXXVeLrnBJ4ik+p7
56RyX0GCAHVed3Tm9kMlqn3oGBI32maDcpSQ7EYXEA5y8ta3TPut3dn5hYsdhsWYlxncQIz2WmWq
oBR+Q6YSDR8XwxeE7d5Tx35Q+5ik8IHdnIXI0AYIPQ+sgGSDq/C6+IeGTrf3WLGQG46dQmoVJvRJ
xAuRcXMRZClFohseYUprveb9JnIF/yvnf8H8gJbPM1OGh7dZaM9ZG1YADxj0vClK8zW4wMXvdQws
+lwIgvBRQ3lnkhVkPF/7911HTVC5pGTlSnEE/Gdhhn29HV11Jke8Xfse1o044pXijL9nByWSAIRD
reXpU1mRc6FxKb0+HUB+TQ1k4ZhkuWlh8LZB3JjUGrEX4pMKc6e+x28QqC9gCui9bRZBXW8Xqa79
O99WyjcoqZzNFtjAfxKH0WkLvptPX9u5dOvfUp9fohrrfjOPUhOlxlMmQuR37L5HZIsnrPU7LLS5
XKke78RcFOXI2hFk4p7xNFpicPkPbgCzzDlfiBXmdn+SxivNgla4Y1eKdWZud87hRRDArPLxVFjq
rK4rbbePTD2/yarPB1m0hjYdP4jc6noLa/Nm2ObW388FpE+jYD4DPX+vVnxPAwet9dpWfP5wCNQb
6CvC1tkrUahN4D32Eb7AonbzSUpCIwLRAr9vRuPVzaeCICqkn+5dzLDTy2Ar4Za3ENbwT9/a0hGU
pULNpfmkg1IU+C++PGk8+He6t2DbHJsS7ucptFsOM0BrxF0i+ADZ7S2YhQBLloVR5gNJ0X9JEkpy
faHzFsCBBHfv03aQVCauNem9GnxZmrZP70oZEdLh+fgRtcDqVir7PMBexiltYe59qYswyPQ3GwGO
cjp6nnvWkZWhKwHYAS3uqpHFqks1p7D+JybmRe0tNs7apb5OsZJBDvqjCnGTkGQI9SWyK3joXGmi
/gDD9gVPhv+fE0j5cfjIzpPJvSvTiCIiA1MIoaa1aYvfcpiH5p36J3Ki+sE70t22lk2bRsmd+njz
/uqxMjX9AIqEUnybv4oNISmdRvwjHsWrsD62ZuHpXavWZEATJtW455hRiXD8lISOiL8y5xnsCV3C
LaMKkKW3+vxPhPQOO5m8mp9+IHSJ7DnYac5VfowIloFZZGVgsuotChBjUrirQLK2OfvaflcHyTzu
cVggEZhjeK+5HKxGAT3Cm5CLoP10c54hRXFFzpLpoPG4rtAhicC4+1eRWBIfjWwZqD5HEoGhsiur
yXga2WtA+2J3dokLYGVJ4B5wASwUEA9kRziw4l7w7VutGrW06mTGG997zYksba0WOx1a/92GK5dD
xrDBUt3dhf+YDig9t8x00JUrQj8A4p2x2x++84fRQ/ae5X63jOMx1ZjmEesG/bdIBgDW6c9yfNhH
7/Rw7HCDNK7e++REyaDyjGzdx52LV6tmw2mbkHmQE09VSeg2WXdgG7B4PtqxksDdu7bwCSvKdKdw
rkQ91P5C4gmLtODxiBlrZ52U5Pzn2/TiYPghI7cJ1Ly1vltpz94I48qiNPNtRShVPJNLPsoaCYwp
eslPo4AL9a59E5/5aThcbbZpO3ozP9u1zr2UF25auup2InE9+Hn9g5EHvd5IIZF7It1/x9iYmGtY
obg0ArqpZi0fbrt+bKuy2lBs59pYJufwXyLso+m1bopgxcQ4bhHxFHLf7DJ+6pMJg/mMXvBElCjr
XySnaVFdyE+AsxfYwknyLyBR/pgiLhxSw+Uo4NvLUY2ftV2rgoIyQEVPQH0NY/qQ/C/5VD7eQLbj
PA9PxTgfWkR6hTnRKWDt1jNQfiBmOd2c5dnWJ0SVX++NlLNCV/PCdjkMYalP5aYJEDL9xnSB1bSf
UQUB3ay/1slH6LXh7oKtLpYLrNsYt0Kj0nEUAPk2IlP1bmtcB4CZOaBxZ3dpGSrvHZxL9fuBxPZJ
ctXBxOUvw9ivht91r9C9zeBc2Gcz6csva+89f+P7JuxjHLgna1PeH9wHPDUe3zO+xqelgtyLj8uW
7f81HieoLY8sH9bFSYB2NBphCRah/6h4kWY7VJ1uUUHuxsmVoX5fl69mzDscee4e8EIeKya/ju2t
yvuUBedd+CtmVItvYdVLiOEgnYRhFrCQMVN3+stUVUuu4lHcrmrU17rF1HOnBuUElV7wRskTqjJ5
/LXY5gVgnXV5QnnbTm0ST6MQi04LIgR1KXsO4ImwsGreLe3I1+i1odsfjLj0r6hiO/fKw1tepF2P
nbIzzLj7diEBsqixWg4RvpqbIFQK/MWNWff1L86JRbOq4G6fVA1Lal4gsqW5crtM/NKkjYvsCB1O
zH2yQUHo6F8m0iF+LKhK/i0D8aiUV7g1Vk7hnEH4nm/Vb9+FN5lhpGbYxJpuQ2Shai6cz/OBF+v/
Nh0JJ4E/CJhKVne8bL0tlUrEzohEgFF82SGBm00xk8KYloTx/2muxocyiebCFEIV4wmfo+RHUlAi
5l2tW0XuqN6ZW/SDyGdSuhlj1tbkYYx2jJyNkNifQa8MSFPc8VlL0694atztO7SxTLYlHLbQ2W37
D552dBUtWDtG5jMfZj9xYwUFjvaeGXziIoGA7Vr+0XwVutSnefJklCyOV0u4d5pRhpM8vUfcj3Cu
6f0xxQ0CYnSLdcp7GJn9gAiGHXOMDHfGr2ELvNiWmURe709WM4w0ASbN49cs7AuCwnnOjIRWi7FF
ANA4PpXI9a2gE3ko2sKbxIeo4vcHZYJCYi33eSiA8AV8U0c1nmR8r9cMKa0pfc7XlcDsavy3bGcA
iZRXzmWRV04muXMShUDJDRYd2eUjxMetTpiunjGcHs0tVkFI51hqDRq/lTPu7s3QENfREuiHHOqM
YhicSEjlbEUX5Z0f1HaqVco47DS3t7ZgXJHP8ozP0XmIOorM2i0fu0/v0ot87DpFccgP6fmoN1n7
BkHHUWjN1D2569XBkPdLFpKNxlTsq9maLBSvRise4YuuUfralGWUTkwXNj/BUouRgDQa3fDfF+Zr
0msWFcqjNV/aBE1Jh9FNz6HIkd44RrDc1Z6nByTbZBDKeSpJAyyCjvD536EQtDUK427pUyjWlBpT
mN9gSLS8gusUTeUGel1h5pre+df6pUZyHHDwRFYaEVydhuXY6NY5VSDxETfAQrbuR3iQtERBrCwO
tuBDcOYRvonwgWG1+sqF+L2wYtR4YrNBPZqWFZS37pt22bVxf0mcJdxQLzpvu35zjcAeQCQr1UFu
xoHl0ptL7j35qY9ps66KJCI/HVTRrTtdSiffEATfRFDp9ZEBQbiEfWCntTcnbIB57Hx7umwnhPBM
Qx3vuHRsE6lrbopdtEaw7UC/iYPGEzWD7tWe5sBdvIf1Nca3QlveNPx7hBl51Tt2PSL7dO0kfew5
dXbRKZeQbY+Lve89jgf2RP0WQNEg6zAqTw2xJeRGDMlDiwubqpbdv/egLqtTNDGMeDfiZMu2f0DF
cyWkA4pN1azzWYZg0KSuZM7jkgsbEQOhs4Iw4bLbnO7CjVbhf0SwUE/RRwabqOTtR/+sFbtb1pY5
yLj3z+VLUmuwOopTNXaLP9Ljf3PbAwXAlzr2zVZre4XOYyrfavoCCR4563dF+Cp9b1U3C60AxAYW
k1SKMxsaawUHGkeLqpSLYN8vUYArhNdRGEHFeesp+d2rKAQSkjNxyNG2fPwQAcxqNWeo2T8jL8w8
jRFaNcJg2xuWkgWnEOgO0u3hDTMH6FFpzV1V394zCM+lqUWWkQd0F2/zsabzjZ9TyTLwEwQrzRwv
oJ4S3Zt+JbjsWzm+jXsE6LtdxNG2ADwfJ+xjbCZjEQQoxV3O5d03+d0jlEDXO7rQPwcpLvpWFCk4
l6GdbahxzceG9/q76TjJGrz96o13mGQQUPatxcDHea01dJ6NkU5zCdNLDO/PRTd0cyRaMYQMF5UR
hBOxXJlIQdSiJsNixrXXkgcaSybDhJaod3ktdpye4DoCXAlanDdL3gr5btwI0cMmHYlvKyo9pAXD
8pLkTR5TwkRlREej2gnKctYA97dxByRuwazsSrfX5OevsITXXTyY3zWO5GSmsRZscEB/JFs5Y9Xu
8nF3bKQzOAo167NRyBKQG37N6Qir1HKS80L4MTS4a3VJeUwnMV9aCJUEGaCuwNPsfavW66E+lKE1
/50Hm4iWARU4cWNJP9sebiPhn0Axem8y2TQYhILgf6C6c+rEYDJ9/fGl9OaBEQL20hUsUiFl/ywK
y9ESCw9lOIejV6H45Xcz+ZCD6URyCO+qq1tFnmAN7WhQw6Cng4tLDZr6LhCMMESNTBDZaFkHnvS7
vBEfV4D/mXxa1Q25WYKH1vl1FRtrb9s2DG8BGZq2m3x+phkFU0ChG6S14geJPX/e4b2Z6df3hkaF
vFdliivV6lgUB0stpffa5q4rxm27je4k48xD+8+fnB5cCS9nqxo2koVbpXsDydz39RR6Ggpl+L2c
2BE9i58ml1RXz0BW6frcCGfgP6/2sfSO6/fTJhZYUVuUNd9vmG3PCO2rFAOYd45EJiwW1BHT9pf+
9YD0WLHll1b7tSEtdThGup1zJk8s4lsAe072uxwTHESUAuB0dMlulFpf6eAGggqA0H26bjZl+IU/
DDS36WqAO2YzytmWazz1MgSy5XMLhIZR/3GQvJohtj+7SWFeR74SoldFkzjt3napST9nVK+1buti
2esEMO2OZyEGQkCun6Y1rk/PxkipIM1HK7qMVsYiezCCSxcg6aDlkRN9tGlKQaXyHFV6G/4WxbE5
BjRzlPj0ZSpZXLP4XGAqOaFC/E01z2X1uK1K/H6dX3GSHU7ESmrpSb7eSf5AiPqyKcGVT5ZTigvT
P68g4aFpcC3lMmi0vP9nT+rb/gutx/v4jNjiZxFDMoOrgCVvl5dmLAxIKA3N6PK7wqXKbiRf34qh
7hkrTH87HUNIZFiUoOg4QlBgNXoMjB8taXcs5/iyyck/4VJshVYC+w8WIlxWmOud630F1XqFThGR
Z5y8iovJY1LMUWmuw2F52+N1Yp3IhCpyJV8IqUr4sBf85bLggUM0vTqra3gh5V5ta8xxreSNZJfW
P6cHS23gkRV/ht8Sfblwa19qQvTtSd+WgIQGQZxh4JOoaOW+NWQIQkgveN9suwIUUs4x4x0crgZh
LIgCCBYwN89wnAFTKC09QPkgG3ND7monIxbHHfqRebsnqt2TWZyYL6Er61Bs53iatH4XYJH3ZfwU
IRXmFpWJ/fPHFlHzWLEjv8XkW4chxri6FeN6ACW5rAQ1qMmO9SVmSLJIjJ03G23aeEq9rXKWZlzi
rqps3rTKb9sF945+ggkPsung9AkbkD5ZxkrS4dgPhC+6mJr3Xau7eOy2KkzC2K3/VWbyEJf/P/Ka
ivUOgNdnDT7e1dcDuVP4qAXpu/ispayAWHYgHQGtyXc4klVQcxRIcKFu9nLB4oxg/B/PaQ++EZf6
5z8Zs1AmrDl1cpHrFBUz1c4+0wIwLObM2ndaMEiMkw+HTywtVhrcoJilxBANO3QJNiXzejqIl5UA
aHO+9e2KNNVZ2Fyp9nufRHiMMlepy46feNGhK3eDIYZ8UOmZv32ft0zupXcEnMeYeatbhf4+B1hI
RXXxmsEOvPO1eSue8afVKyeYcZwJfK+Z3XKS5/1v4CwLwh+6RgKczEATwv7MJP5DVT0+NrdY3xrx
umypjvSd2J6GyYsM82ld21YWQKN2kxIdxT7qj7ZIJdhyoV0jMxMFxCM1QqxT/T4AeUtJRwus/fcP
Ru9YXn/fHcmH9AHIHu8xjFuBXuoE5mvFRtnoOfkAp9zV8A/qqistEQHyTIY5wWw5boy2+SRF70E1
zG8QfGyQmIaQ0zwyNNiSO9PjcYtTFl8YF526O52lYM6hxM4ZdtasWR4Ro7sZpKLuj/rqVYnrayef
mLSK/jXjc7MiqCgESp39i4oet6km6EGO/hnGahtN63O6+yrhQEDi/zF79zo2fsdD1KY3c79mqa/K
WQnGz2hFdQrocacG32mEwOnwEmMp6quezkesOxa+mbpYQQPkIshCDA7qLKN08mCuqaLmYRR0uY5V
91BC50+3bhVAWrjE6CCzjS/X62lOGy8jyhjukmIS5Z+BdW24N/IB/7Cwvc/H3XCu8rKbpqPZ0nX7
MPUpplyE0IoggSy3FSJNBDIEyxIcQUA0XIbSiu0UHfiCGjFL8Uu9wUhp2k/nwNDQEbqzBam594yn
uN5sZabPzUnE+QvQ9ijp0+dCFsrxYntSF4nXxwTyZQjW9Vnt/y/sXZz8kNrOqRwFvnoqvVcPaJkl
FXIvekXN7qTzmDRITi2Njnyj2SED2AoKI2IlkoNfeVjgZSp7LndDyxa1kqgyQ+Z5sfqNvOym8mrt
qIfs0HT5EYlXJm8+L+QFG0WEaj2yp/L9LYMATBs02cnQgqonmQjexl5SfEJNIcFkHDGfUWbLQlHw
eWUB+/Hgc7fJXkjXDzwqCWownatUhc5+z3xYnhsknRHiC2wlz9+5gVZhoQ6hvNhaHsN/r7iLA3CO
iSibtjRUFDtO7nrl1wC6emLTYHcVRWIXCVLl3rHcee1pT5zcDCRD1797NEfRXz+6RR8dj7Cz7gib
CDJ6BSZXA10xZ38yiFaC83CYMzKRLm0vBGcUhIjxrQ7+7mEX3+lstnO/8WVWUREUIqZvgKZEkOx/
I/eo6QVkTiCpzTmw7B0csm9tHqq/QOTK7diPvTeeLALU+DJ3hKOdQHDCqxtXlsrEU5e36uZTTjUN
sDHnctevhekeZfAaQkLBSzxjUAM1Xbhwr7plgXOINcDBiEl+mUjqf+QYDTM2KQ6tlemjsmLpHNDN
Tea0Dmx4mq4EGfiv1qNIDJ19HG9441uuG0Y0p2aGvXrnh8AAG9/CwkPpTRvIwOjzBDbvMo7Rwp9J
NB/bXjqbw2ox7Itq+MAuSk3uQRvuITsvyaPZlcoUi0oPoqNwOU3FbdK8UaktVHHLFPO5IMB1UOQf
uewdUyxWD6C+wsl7fYPHTfxf5dmsOfPGuOdq8h3BpJNBAcAdBqPs6HtTaqbk7pBXlgbms1wSpd5G
NtQzZ2UGJsrXRe0GmTN1bxr4B1mtS/mkp9TfEUMGOUz7al9VBhvOnRLsJcRkC4zBAwO19O6+94+L
KJWzwPPkYx2JHuHjp39cAHCVfXCfr14B1Ab+6bC3OH9WOPsZFzm/UHmTVtuWUqi9PnSk3To5uuh/
bSc68t3hVaM80UInFHMh2YL8PD5HR3ewrT/b7CEau8F4IINaT7912bsdDUZ+YQzF5a8EVAiC0MNg
55pWwSYciyAKEx9eTqplcBwWsce3f75sh1Gjr7TEtID6TTny3gwkomtERRoi2628+wKYVj51gJyk
kdtO4Gx0O4luJr7GlyJaX5kbJSl8S17vF/ywhNC0rPRn/Mu8geB+yIKJLsdpWUVhAueSKKYD6NCr
8p13Smez+0OQGPpXHkyFhwMPwSVNS3yvn8G+vKNr19eb7g7/cffagQ+O8A6wRXUIa0LI3WdOmJoV
cHy1H7cLfp4Rw1COKesEv9GI9QZDo7Fn14d39xjGTE3bwx9j24BVPY8RR4sD+mBYvG4Lju6dbgdn
RQQsDitTQKfeZ41Ov5ZZXWKqyvCjeIu4mFjIublykvRuhpa3P4GP6H6yd5nbagI3YIUMGpUnKkPi
0XSw/9OGt4PGYhm10eeCmbx2eksU+jIp5WGlb/3EYcYNeuAHbXrDYlE8GTtJ2v9gAuvRnyXaYl8p
0Tx2/lJJ9sI0DdIU443fg9/7oNS2J3Dztn7lfaS15AC20M8/69Pw+jT3Pa2kfW4UVqVAf5pdtyJ7
Kp9gwXFgggdXhLbPU48qQkVCcDhUzyMM2UYKK3R8EpQEhBOE8blL4MYStPW53/3m2mRcByN3veGB
Qf90r6cYoTNwmxUNH/hXKxaRP+ww1XnTmmmmd39le59mqf8w/n3cbzmD5d87et2HKXmSidIP1qKf
qcS9/AoKIKElGtvQ6zkHmy5Aibts0OuvaYYZoE9mosewNg7IAqeJOf1d3VgrbSog7rhZHbWgqXTM
HR3Sno/unUPvSTycFr1zJ3mvkhwTNH0+sX8ZCTkFy33br14hJPsik1qCrvo6cSRtRz9XxNgKBpOM
XIzzxOjpu0TDw7/zkFQgycW3HRH8fWcrjW3B3B3bcMO/n8MB/YwbxY9da6xGpOEO2pcu/EQKdZaW
SY0kxtIUwweNnE+mistswwETifGyhxs/XyPrz3gLzBYl33S77temQBW66I4LRTuvy2y9l+1rEU4n
uM2qRRi4lU5l6xhR+g4UQ1SowascWhbg3xVl3+fprQJSxe7k/0EXpLFSJIZro9aF7BcCb+CzZO45
0NZlHwR6J3JMDxTZai/K+ZR+bfmdZVawm8wS8Hx20tyvX9+Moc12/h0B+9MhfOKxWtYSan2nIJgJ
g1skiDj3QMS8JGKcx2GJYlACTpJevBHYizioGuawvZn2xN1pQzaqjPFSXKy/CyyEqpeu5yQlXNZI
SDCWKeiN13M4D/wQZ682xlEXyaP0FQJvsBTHn04px7Ly82WH7bph6N0TCrbLHDPFOVVNjpxCGlz8
b544pb3iq867KYaIKbarqG+DHs47a25D97j2r3ejTmZGmMnOo4MKxvn6oxifA3vQthUlCoTWA25v
zYIAw9xwEiFZ2Kuhp/VHJ7DhRrJrOBxdUQelFYQWc4pANqU3yBxWY3mrEkn4aU2pRc17eN/kxrbp
d8dBBQF/wueryd4zbzxI4nuTIQKLwgkR4Z1k64MCJPozmpGRGyiLR7wAGhIWRuGFCDL3Mp8i0nNo
z+CXGiAZG8c8p9wkaKAUuuKuVGnnI5H89MmYBx1vfo3ppB2MV//4vlUHA+toEAxfEajycZ38rtrX
AIpX0cIYEOns8rkQp/Wj7EE0SMz2gX6R6Pf8e1pBHUq1iPXPgrMfMWTln5JyYwHgiwwmBKDeHv9x
7l5/6iDEWvEJ8fa3/ktIsTX/rbp5pAYZ6zHxCOO5r6UBbL0fWQjhqm807pLzbYF6kYhOwCa0nXd4
LxvLGA2L8Yqp1QRCSW1+ueoGTrtAgdQ0bsGMxw8YtPGfewL6yKKN3lKSL9MEQ2oYjXmSGiu8i5IG
CNtlUvYtvEvbaxDypUSS9mews72fE3KlVLfyHgNiiILMq3liOS7Q/UNfLELqaRTZB8cT8/m24Zxf
n23WK8CNZjIyIok/jMrmg2c+CXRHydJ4gMhqSGD8cpW0jab+sSD86av0h/PW7KTi1sQuntqTodNC
AeR8dn5G75A79Gtg9yIZn/1JZ2lCI2WBOUc6Ags7THuF8eD27WHHONEzGex/9Vbb7E9m/7JQUeoY
DUpFxBSkKe2KyaTXSAgN76Zpm74DRl8tWfElMVKqylC++8HFbYOBRZLOAmkWIBkBevvym7DfRgDv
CqtnddRubWmrNaSHo5u9GLx7yh9v2doiBNBGYrQQOx0PePVYlvoEcrV6PFXmBNVMUHPLyiPkTqec
8r18Db2CIIymV/pkO5mTIZ4t83eUQCq2lOEljfQZ2HBs9J6DF+swIO+74qpSkSM+pQhi7PIDXwIq
Ho7EwENGEuf8LhF2s/PV5oPXiLuoPUcD5m9akAP0hmgnmsGAxCPJ8vqp9SrU4iT6+GzqrIRVcMCB
I7VDuFAnJjYlQiN5b2ljqMa+9ZyMc75YV+gs5SDIhAWLKtk2qzII7pvnStw6uYwFEzqQnXXBYg+G
g8XbOdZ6gagk/TpKKyH0k/hdf/1Hy5hj0gwWDNJX1TnlwNbpfOfYjt/yDHO8tF2k4y9KTshkwdl/
UGuRbyz2pvVv3/Bo57oACBOvu8n271CI4Fz3AmU+kT6rcHnvHazWYS9HPl0MrWS3ZMTE5PZfZZ1O
x2oNP/fXljtG1IJ+Vd60uU8XRUcbPPsk0RgD/QlX1Qdv7Y4jRt4kCu+ZNhKBW8IvRCvBdKIXWSx/
lEP2TWyG1a8g6bIWGb8zqLeThSeBNnI9iM7uC9uP8YBdETM15uJ97fBlzjfObG7FsKkoVnPyLA3Q
KcDKdGzM0QhUwSiYHLdG3dfIQIkdNycriowva6jpZTUrCARP/9wr3BamtDsCS+kK35HJ1TwgS163
WdVr5li/jCEwXn6TuwZrBIoY0bMTitOkuLbjLSkDSz1yGr18z5mKhjhHL8JQF+2Ea3Yl4XcZ/Oox
z3e7FKJAMuTFga6Ho8IuSv/Pv1HsBnzCucqN/VDOqnjmZuIxtOjXMbx6AmofVR4PuhwRg1xM0mr5
5Lw0xSyZ/CQF8S0ajvImnMQLJcsVKSetakFAnL0a88yPPDoBgYzRlaoJ4VJpLxvV/zlVV1INHOo5
zhQ4UnCvWAE/Av4yQ3/FnKT1Go2QFigwm8pH9yYOcxk/t3TxJTo671lRoJkQIIGX+xilsYJRiuPk
TSFotXa3bFtdiNJ+UIO4qytieeVIe/QLf7Vacna5MdJCH/a+5LSidDdznxdg9HMk3pklSrUTrp4K
TqAyVO5n6qkrpcRxQOG9FP6CP6Y4H2LKi9YQa1D0RIUCTZPTG/uIGG86nKeMe3jEPt81BoPkdui1
uC3acPObKTD5qUUF568uOorQoeSDjs1g5P5Yw9tt85UX10CsRgssKV2XR7UJKc5EyABZ3k2htk2N
RU97p4dUaQh4lOEbkI9dPMgWZEnBWCtwxo/TXIEsqlAnm/dBhPyi0Qit2Dmczi/49+u08Np0M86A
Q8ZYdnhCbIsvUYVE7hCVvYpjjE3DH3nTxdL9cUFsEBYaTjakmCbYg1vQHd1uq2GMTj9jewbIvXdN
88DpCsPN61kKD40b/r1FPRUzKA62xH5gbpVfJ1eAidOdai3rdWDRiif0oBSi3k6ZQovyncR00vAW
rL+4GssxvXUUvDZ/RrcpBqFZb4HqQQnk+IjwXkpS8mtqDDg75KAz+XUP0gUnSkCgNp8/xn4yKc1j
gV4CLJAEIKo84sK5BCVpaZ/yM9rco2JEm6VrhuxhQ8pIdftcZnfCYcDkEik7jn6FuDyFEC1kJ0d7
sgzsfZfxass6Sz6ny+EjJYN1lxmOOqqyFoMAILRypl23NCdHR1mZFrRIbqKt6GnRrUqyrF/wcrdB
nte7b4MG4apThya3u3dS0/VQg2Fh/OONMKtutSOf8uTyAzpQ6Mih7qyVzuy6tQz/EjcsOCqe1dk9
/BqZKn1BojhIpghUM2XCiUfMM2NEfg7iLqjv8UAv49QTTAvkCGN/yk0P19KJYVGCbt9iKTjFlzq3
uU+rUq7pAqTyhXYz06dvOw4AxZna4A/1Rxu+zZWUhfQ9u5QHnn1fKj02Uoe3Es7HTG7INBQ8gXli
UaRk7ngQj04HzGSbpHwec2vdsqK+4M4mFInMniWCJrlE6/0EenSBfcxccI5kuHMACk5thkavwMla
xfQybwK307lyyHJNfDujRtH84JscdhB0VuqmFrFrzJWxHGlOh8mr6a80PXKbDwMPl1+cxYXg1HFS
0mEhA6qC6VWHEoqcz0tVNIJ0K0NjAaPCKxw9Zdak/x1eUqwrgcf1St1xzjbrpwXom/XYM1deLMqB
DXOCOF7VTiFNJiRijuRXE/zHQL8WhKiERHvtY54hIsw9po33bvgYRbgzlRM19jV3uC0Nq0UMy24q
/tLeFvJi0Ns5gXTXteeSjBN22VuN1g4yeUlQKn9HL3dAbWQpQ8uvzN6FfrCZsvBZa9wkYFKrPb3e
RbYbZgyQrHAja5uXTbehV68x3ZGMiCCyeQCYmRooJTLCnblTw6JLZfI1xF/F/3uMt4l2gk1RBSUE
DJs8JUFrHfLTS6BegDtRZ4kY4LOl5yHg6MBvH/aiJej/04tQYgXwMqnKS3rj00f0GHxlrOH3k2oP
HtQ83Q1NkZvneujyqrkZB7/ISsruPylkkZKAnbOD3OaoH3Br8o4PgqLudk6+7HgtteLai/yhXIkH
3Y3uKHot4LJ7ODavHmZkBh9sSxAIbnUDVak+7iSeEuQStI6JntF8MxqX+6Q5RpfLjddbr0jO1Q96
/PAWRNgH4jUFWyGWiIn970ET4ivnvyj4rtj9sroWXTFYX6mDDIbAnvJli4Q4tcXzcuvh4+YFZnKa
uYKwXzmOzIdZO3q8iwLRCWo2krm1fYyQ7QY68emcdgfcUaw/p0oa8d0I6X6BnsFC3FxbN7dOPdJM
qschPDWAlkSrmYodhQH6IY5+SexRK3+becGgUpns0T992RKM/PMES2LHpEbX8NoNX3hJ6qqKgHlQ
cG6eLwyIYdP2kbAqm2WKvh8YhwzlmKpAaphDlO4WUKGWbjuF7OP8fsSdt4kqM4ypfQjMMX6GiSg0
YGCLibEht7JX5aM7IGv3kc5qmQCF/EYO2hxjaLGyREsMrUgbsNrYEBTys0Gy28OZxBVqGPwRHi3I
/h00e6sWP/zLnEeRiUyuHqnUiSAJhE7bCWYADxG4EGMs6V+XSvo6PEi2K8Gxf8yH0PD0k1kwjC+d
BKatBKLr7I8PJc/qKclI40LLX1JspQGjzwHwiozkSJN48WX13Z2k360sswvizHYbcd7BqFof5Rpn
LYzIK7X/s2KLK7m+iy3t+iH7VLPmrwUmYQTpUFjUcRKs2FDoqtxephhF1gFwfaasbSr8u2ueJogM
nAbNzQs1MYyWwfUU69wicXk44nPyOuU5Ydf4ekXeclkdmsuzl5logpR4baA7+1gHnX5n7OQ7n7/J
0fSmPZZLjOAMb3hF12EUhHJeNMbLwx/LGmhnxZDqPkGMCkm7BO7f67YUFxZAGD0fpuK66/jU8kZD
tHU/Un0kJ7ky5gd3jItkCN1rRnxVDqNcMszWNy2otxm/huLDA8p+OVzgBLNYonr2vNhLSOVF4plX
aWDl4kM2D2nR+4qZpYHeX1DwnAPNPC5IyY8Jho29ngfR6+QzKXJrpiszKLHCbyVrt21TWEW+J0C/
CKgQcVV1bo63WXrkbVJBne7DcpQ/4dQqfaFmOYuiYtYlA3+rZpbreTYzlEiuN/FsBzzymyn71D5k
8BEDbs1NlPfzuQpabr8Lv8RMe2lMVs9OWRfs0k/QdbEUFZGnTAfU9KyCpYEqA4PU4rEcqiPuh+ZF
XZRZKuJNzO90WtGAMJCnpB+7lOyywzysbmyf8l9uoeT+m4ug4IBkM+6snqNybBEZJU7yQGHfOdK2
FM2K/bOhLJEH5hRLTVDEFVb6v/hP1ZDLR+FaRQv2DfQwMLP09saNUYCRtG7CW+9mpfbDSTBX3nUu
j4iovSNc6wxGO1gIWGI1NDZIZaooDGYq9Mc8j6F/OJss0RM+c8zHlHfTejED9oIQBzUA/eW0LUXE
Ds84UDwYBoUCidhxoF6P9bNi6Go4hQDfa2DjMDKFrxGwYseddHSKmIE9OtaARy5G4VlrclKSVH53
dp7AMNop9KEkX4AxzHg5qZ/WbaF17qXGuYUgGzNGV//l2d566b2DFOqPTU8sf62+rB+K0I2DvcHR
A5r4wbboAEmCx9JYwam85AvDsVmigpMJ4bm2hdQ8hix82Ewxpsa4nm4i5IGdfDI1Al0MAHpu8vtG
62/PP5qdYhU8lOAR6JphhPYMAtJUcYNiyeuD7THHWrkuienXEKKBDI9KD+00hXY50KEPval/Homv
47yu/RsFwb6+TUce5zTTVq940ZzNgWDiXQ4TkMkOH8og3GeZWm1TpUH7yMGStrcfvgp0hyA+Cupl
wvZaeQJ2ttoz7LGvmYcsDFiqmcTIdXKmr1gbdOvCsXHM7zoYzbBvalX6sRYAuU9N0FwEwKe2LZQu
4GauNTxT8yKoPqSGHduI2DfYzpiNaDCbOGXoB0eguh9uFZKUI5h1X9BlbFC9UOnwc6tfIOy4KnYY
Ss4V/d6W2Ic5xhalZ2085Iro5Nj8WP7N3VsGJozmwOYVaPuhjCw2ooiWFSPTMSTfPPFw33shWm90
zn5iyU2f47F5IcjQt0iftGnA1AJISIozPxEwyIUrW8ssb90glR7iykJJ2iVUikgCqWzF568fIJ/p
0aJWUdG3d+Zs6PT8jzngYKZ+0TkccUmjtfe4SHhPpjBS7JrZirfmI/Jb8bXg8Ki98KpPVilKv89J
mUrx5oBVaY/FGINN2ClA6GXaH2UH19BfItTkHIY2bi8BWjWYRflfrmP9JGIlSEum40u5ggrQr0wS
cqcUSGtoCOserv78KLrvLQRiRp3OySO7xKfObyA+ikTQCh8VSc0/OwKgjBuhDLq0wQdHuq24rt1t
Lmcz6dbBpH9t3h6AxjRO+NPXmEPYvYzfko7JNiWubCTGeZfqKA8V8Yyi36+sXfraITuEs4UKimMJ
o7isGuoxXW79oXcTmzffQlRH1q6VqIuzkgTasWUVH9uAh2GYbur7xZMSHk9NeVPwOOIfPCuPaIgj
aPPJ1bDGezr45VXgAAwOIabyxLw+n1MYVd11X0H21mckori89jDSj6mKJxrPOQQlqBewI05acv1k
pVFzAtdIaa17n+uvxfQIy6xSfAtGUsQWnduRWI0K+7Awp7Ac1KSOfpXoZLdwwbORU/Sm0OUGASaT
uYjCjZoCEjcZh5jrZmrMv1MJ3OJELTXuQe8XT4czr65KTQ6kN1csut+n3a9dE3VKegefjq7pG/DA
0g7rOw0F4hAzsbDGyEzim3LETiRXpNxivsg3DJu5+cMQseH+AvFl76ale/PijvXo7I9H1JzR4mrg
BjlEgWWuDIHMWthsCESaH+J3CqsCqe0BA2iq3GcC6TmJ+P8My+v55v+R6HIRlCb+Ye2gaomLS1VG
77/VxbTr5Btxo4V1en/bLOt7tnZhc5lpB7eMZS3MI8XR69sAlkm8b1a/Echg4S8u/gd6BszhEs3Z
HwRzQalZb1vndncByW8uOKYGP5ttARPaW2NFghJP5WNILT6DOHJwiIDXHRxLJIKvtqxlgA/NyJnx
NkFYsm/JckrxQbVMHcfyHFqasX38g20mBZTKiOfN2b+afctrIem1hbl49112Uo1kxhnC5yfhr/CY
hbPRrF3LFZsH1NkLQzat+ipvYil1XkWNAIPgF96ixl3c/X3HTF/+g7ZRqEs5zo1CHiFhMvdU0Lrv
+yE4IKYOT+8fQhkDqudLkK+Rmiif6ESXTSCkTaVM763yBrOAoojE2wf5ufsZ85tTNwAmyMD9Ngno
fHrOihQb2uMUeoweMiKwfaUZ5+1wdrL0iYs7NfPJos7RnjYDVSWWKikqd8wK24pTDBKN/QDdSfD8
tpA3trfgdAlcs8PjfNblFviRghnKJEvVHBgYeAOXUFHfpgi68Db5aziKBRCPH65lCCzJNSSY9UQa
xjt0KA5r5lNrznNKwE2vLNZkz2tFl84cpi/UovQ/cpL0lt9tL9dOg+VNlwWCaHGvI9mrGT8NWrKw
jun6qxg5vEXg3K0amaYZ/CMYK5R7STUyBBYazRwb2J9ur3UcerL4M/Xmm0B0em8RM7G39qcu7aBs
Jyrdr4BeOXe/lM8aAx1LXCnqihSGGVuPUmpNbRfz3uReghh3F6mOGKUkP31oEvgetNXw3xM1RDH8
SWqjgMEgGO77Shr0xPo7c1oFi8laGcY2Krmm09BapfL3jM1kMF6jVAPFMliMpjLbN+ruXeJTrznb
HF/WPmrTPwT6ZRvkL6OVf9TZRbe+80j4rKrbO2BSVaYJzoxn/J7rk7QxNXzstOGqqOM3ARqmpbL0
RF/CzANBtzj3OdSITum3w8OM/rVDZo15ruAddoGcRnLkJoidQYYHyZFVDKlZ7XDRc09QSIRpVpIT
GsUajPc9qSeyRf7KCSkIJi8CZqcjk47oJ/iqADp3rVbH5TkYewlrc2SFt9FmFOAg/EpL2p4ABQmu
Y25sEIrOGmzVwFYm4/xJMDZsOmJajMPoGkWqGNQtN/YbuWJ75jmMeCMDdq1T+arpw8fWZyKQhmpY
ZqkdvfDfIVVDyBGWPbzU/yCON3n8BFqKLRGZ48khL5MjcQC1CklxxZcsfdRiVnL+XfyDUfHr0JYl
m7gFS5NRs4REDhyeHnNtt835jZRUM+Fa3TC32v0gJbxT3QzkjNkPVosJ5M5b6F6chD8ycDCJmGZc
JJkji/ZtT69H/3AA5NcGC5UPKLlHxLqG5eKqX/8e1FB4sJ93GSzplrlxIt6tQjol3eDJ1YrQkder
waDTS3bf6S2qRZ9fuAovhsf24IFprm0HJB2DO04ebmUJwF7yl57POnc0OwxuPaxJ9Bnx41ROyYBh
fnrYRDzC88yxIZU4aew1q8ukZXCiJOg736+uai4WuXJRGhfOPQSLc2PHTDzhILz7tZIzKVu4B293
fNeYmEVnBNrZfSrhoeRaSBzExkNitG6i//uEFbWVWwp9cIbDtDUFhrF9RjwpnyPcffS5jknCUQXK
ekEL0dpVa1TFi9h87LwbwWmm5Cy+MQdNQJUFEbPmlc7/q+csPo+taGplI1/ZuU3soXEUo9hDi1ER
iM4tfMqknKOuK8aT+9XVjV9jAJ2RekN/hBgpcvQP4ykYQgr3H8zbQbIiguKKaR5XTTgpvQ3RuXhK
gUunKw1UaDdxbi7bAemJrdJmANdvbuxVdsFJNvpCJC/gdVbPJKTyLyWteG4g2RLf2wSxIMySn+nX
WYzkiB46vKKJEVoHXGPF0H8TlywTcNwoLekVop03kw2BSp/z0r6PepmCiHS0GavCNCKIZhqh3Xgw
8bWZi65lbZYsPzjuQJVoe/3EeBeCBPhlsLZ6K21syQYTUJs3CxkhYpHUjzskdBvSFbbixvIIsvrG
ljHLRkpQAvBMaxnvdEEY4THIhAfVmTTS6gKYcUmKm0knZbTvH5ktqxcVB4Fg5bgWWiBCZVWXnfT3
kNter7jx/BfLOzV7OFHjtujdOiQhnDQwi9aE0MRagKuljO1VbzVMrv1hLs7EnHEX2fF0+07spZx7
qTJ1oY2IuADjHK+lJXJpdG0uHYnC7Krs54QnITfPJgZQboZHfUMvkcy+d2/nQms5kA7i14sLFqkx
cTKWLCvuCQWJRetwCLttkGHpNyXaJ/8E+vQ6CpYR9IiDVTEd3AtqN9gawzhWzn9DxzZZVVIYUBzy
h/PN57+hwZ4o0W2AMfBGA1ZWxVDecChOMEk502UVe3rbOf1cfa33vXtf66FARqIEdnF/lQlenDIb
9B7hTkK4S1nBUsJw6GvvXsUEfbWvbygJOg/OwVe8oaN/Va7ehXkBzLycBynpew1UcX2WBbIR9eO1
Oz4fg/NKCm23JfOw/Iq3OJVQgzty0i0l/99ndzVYuHEEFMj8cB1qeuGVIkcfznHvxBG/Ls9Jpu1S
RS0NRdt04myYeiGVdc212lX+O98lRtZ/e/566igyTqP8GmVxUbdM7stMZNvP6jDQciToLzy14RBM
0/N4XP9s1rDsNiXq07Fuz6VdMQLMqkYVzy073pPj2DzU23pXxqF8C4djM52CU5UtTyZg9epMy7rf
YWuVx83tyRvv5OxfdpW6tQApmNbFuMfyZy02diHDNlqaa5TO58E0K+9g64gVMvfdsuty/MPgBUx+
bVIoItlyxUdEJ8MjyUMS/KllatzxjaDBv2ooCdemDXkni+vbjYTPuaFCf3XHsf5DMqp0pYvcAuT9
3pHAMCFwZr1wtdpRxGYFScXJN1FZGq2QtiXGKBXCBv355q+76H/lTY8NZnnOOwt8sMjM0JlP9MqA
2TQlCIbKpdFeqX3rU+ZTlJJpGQOBAoRV8emxd9UnehpLAr5cAIZKWuv9bUXpW31XXR5LI+yhdOki
xfS6EfNWRWRYJ2b80AdtmslJj3Op0DfvMXW2dshr0shcnpvaZOZQ//Wc/jmKYSSt8eP2JkLNFf0M
PJPN/ZySn1BWjU507MRz5lq5zgO8j6mk+Zt/F2A+WBq+Manbxo4OLqNEAzXVssjBRp/vNpL3Gcry
B3SYoTizfv68GS5CysCAcGJcRUYFmdFXa5K8gSPhR4pN4l06VU42sz3PFwWLenZ2y72FDqh0p6JU
+aL1dvSQDtlJnHKnwVHFACHbbs/6WbWY+kSLuE/n1QQx//F6m/jJSaMo6r//jMKrIVuYjMExWg8l
a6OkPQtGw2KJkM3AlwESgPOMunXB69Mok/QqeYDzFnBH1mHuJ0U4LcnHyQ27UjNAgRNe2S4vtp99
OFORXPgF4fpIgad6vsvkEcm1YDzMEq7lO7C/kHlElVEGCeNFatWtYoM8QrH8oKSG05WkMdSAJAIf
lc8I6XOEwk+tqXgtPlh4aJQWZbtfaEisHnejV9PlwPXzI9Gfr5nyBz1/cLju3kiPt5PEN9lXckGy
NVtoldELHa3KjVwwzx5Y9zWPq1A1QLu0gb2tP2VIwq8cOnTYeX9fYrQChpj8qhui6Jd5dcWPB4Dz
FFUK0x6CC5RkZY9h19hFrfxFrzusW72eCR+vk2gFVVnPyT+jLJnSb6Wg1X0j4MGhrRciDaxK6Oqx
zalYp7ThUijqO4kX0qlGC4wCUrEL4/IhFAh6qAIgef+W9JQZHQlTb2oDFdXB4JjPDZ0k2JQbQZ4W
Ql8iru+WHQRkDUGjYMwD7QqhQ6G565U/gObicHNUvtWqPjVX6epOtS+t/feWSJhZbejmW41KeXGC
cjTbRqiecEH+Izdcg/GFIiOkJqPltXElNnvOyrRRn2LeSKfjNbS48DM+2/FML6QhBvj/5Zt4nzUb
qbApmUoayW2TZCAvh0GjsKlbDWyO/fE2T6Axgvt3v15LxFULq1G9dt51RtDA5DXUVSebzhfPCBJu
mnoODtTOP4yeL0JesJOtpqBDK5Ej5MrmZneumx/2isQL7Q2co8I72UZn1yymonb/OqhnN2iREVIi
aSvHhbowtp/LiMjg5UYp2wML2PzuBdrGmlxo2wLVY1gzbUGvTqWMC+HzY1B0yQ0pdxvlGEDEJXsY
ScJ/f8t70Wm8eRRCNXYp2nAJ2adsjwD5kYDL6//PEQl9Q5oIO4gZrJ42M3DbNLZakLS0wmha04wE
i03YB6HkPaUC/iEHt4p6pjlPog/ClqJfx/2AsuOLtdC+RuxPIGBQOSwuNAtqGQINEgZbgbl1+vfV
Di5OjNbqP4CvZ/qdJhydDJyy2rvtVpIJDlEp3R6hEdD9LmlwhCKybo9lhAfhbKdGqZqRa9SXW4oM
v3SVu9mSO5v+Za6umv8BWXV8D1Mk2/0iitv20YbHvSeMLvSBgNSggxTqigwZy7qc16NhAt5PvSJE
DZHfobP93hwGIqvpVNdT7rPckSPGvuHs20Cl9Vv78H/P+pB/fTPnIV+3emvDdUj0U8azPabV6t9O
r5DVgi4N2yXsOESg8SAjrEA7UZ3ceZojTwrrKYpEphZCV14UOCJSMVT4dpNbk4WEiAgHvh2JhAea
jwVygvXp0VP329+nHNmC9gxOq4hkkOCttNhSjKwnEpZOaU31lb2y12tzPIwz/xDpL281AXSwjbI4
NQRexoBe5WTkRvj64L7cAQz8OCEZOTIwFLSVN9htByHZlCR3wVnxsyuZE93qR+Yb7FvQkqqCM1V2
kb1gMy5c+eDa8Kgm23XpfznBjWMniFp4AEuPK50Qo5qDOq7M0m6+0df0cX5PbUZHEWT3cj3SJZC7
pCd2sAXusjSXdh48kAy+8L8pzz2Ky+DA6NgtfYV+7glChN2eeL3kOEszEJxLfQu+kRsN3gbpBcbU
DM8Z8RkGbEvvBLGOm7GyTOrHGTmH+B0ibKbgS7ez2Tb7OSybWs5mIWP+jGHpKPOiPXJyz5zya3Oj
1SBwSY482IMixh0KoLlADPBSzJOrYTPE8wKUj/tKRGvV13jesuoMLy7zrW5+Fu0Fe5GdVQA/V2lq
TnKnlqzlqxBSFlcjlyFsmA8YYPpy3FLZXqb+XMtQdp//uPXfizx5rUogOipxy0UmTPsmPNRCSgyI
Ts9vRuWTzsXxrQqj/WPq6arT+kWrX9HHqWSR4ay2LA7FyYN0G3k68Rt185zp4Svq3Lq7d+P/NuB+
tHKq9DCQ1l1o2ckSu1KtrXvrpbku6/V/kU9hOlWeo7l1nVI8WEQTCejW+37icN19iX4IhkXWjHia
cW6cDtjzCCzOmMXbeN3x1ICF/Dbgdk43zVD+mbtztzu+EwGCLT8dFG6w0fE4AqVyThgM7sB1yRZN
xHqeA7Ha9Kc2ToFpFRaXBaxq/c85xcSlY7YuseibI3NeWvxFcvHlR4rWHhTEa7ACWaqgFG4Nku7l
E2gvPPjVz+2hUgR5KauPsWA2JKP76CjA/1kFYwq5m1OsJQy+D9DWieXJAHIWl5q8pWifT2ROzbo+
3LhwGuOQvry9Zd7YyvJsWfFKQRS9vyHkVsYPSqQCvvTxRKw0w3SlzaVAQ4NcCXaG/lRxaKuJXaKb
qi0YdqO3rdQYL0QjyAbFY5kGZrdM7NNG6Gs0X6Dod5p59E+/TIb/KLddynwJeZDy+NL2GqNMLz5c
w4Gq81onjby5Kh0ETh5b7STWmCHOSLJc2GTTAcaYV17dvILOhGHtDcFlqv2HMS1T9AbqjXbACq3h
NEnys6YtPLdJX+KPFClLJKR+hjZoqmf14Yp0OxJGiBIWRt+6Y/3kiYrJ7+Z57G1UyWqX4k0dXWfF
tXr3NE2NqLkULYManFNWwh+U8rrZA26h3YT5wkYMa0HfiRL2AgUX57hoTHsabcrUByrfRs4RQj3f
qc3CShNDbzZmSTl2RaLHJGWEPt0LZE6Ty+RcQ5F6UEOv3X8Npq5+xqK7XK1vvLgVQodPn6BRBKfz
Sq/ZOC6UjPvT7s4Ev5m9iGXXsKSDl5eHSXou8CyNhG9UM0jOcJ7UfRLRVJxpx4jTsIWnGEOQA2Y2
pLtnkfbOoht2kPRSb14I5YuEj5520SyXJtZyH5CuzmAM/UG5n6Bb1SeTrQqWyli11sRnvaDf2rQg
gzpmHPWmpEzIh8pGXcRCTzfIVtugUJj4UpkDRooPvCXkZf+oDw7Fq1VF/dkyxwlHXv5wo7+mzRcP
XD7UcEEbgfHff1Br5H8NExw5T7ch0LmS+YXeuA7Btscc2KOHr47oYA55dxdUasbqyPU6rm+ZF+UQ
0TyyC6Y5prRireymt3Jc1ZeGrIN2wszvJve1GOOSlPgLqcZ1lo7DTLHz+IkgVrOarOWfQO+0/hVQ
IGrRp78s8NXkW23daCadQLMGPagJY9HNY6aSFf8o2pNNqoUaIw7kr35AWfTer75RIKoamKVnLBk/
V1jGLis7up/9gwNauW2PdPGVa3Sg9j5BUp9UGd7Fh4XTTTZh2tabYxzUuwRtE1AIVgWyH8feSf40
8zRF4QvWajPIUvlwgBLeh7kmSypN4dJyLs45Cj+vOqwcC6/sKabCf4F9w2Jw8GBIgPrjV7tQQBV2
izOYD0cUG12ijbQv9VjGz3uzkt0jXj0dJdJs0srlEAgnNAxyAok0smYVOnyhdudhL5JSxQzDOyd+
ePvA2BMEEyGnVkesr4fme6+Fh3UfEvUH3UCspKs3MCqPITnDIyf6nci2loKYwUZ4B9MsTxm3BT7b
iNAGNqF5NP/qm//Js0i5JT3xv5Q5NZ3YrgD9zO4TRo9eGrTAYw5JV6orBkDgXGLV8YMtcUE6VmbQ
3fbNbTxdj0+ckfHkcLg98gDWJXA/PufmTniez1EKjquuHt74v7gWSF3CQ9T3powlBKwCz9fJDHuZ
5Y4rEv6rdUcum4TdWSFlZRdjRwHksYjKwa+PTCoNyGSt2KVGggHeDLGJKi1LGhJGG2qKIROC3ASq
00ZU3eGZI2xfnoJX1TPT/9oK/iRv1mqQ5nW+AtMurFHrKo7TGi+Sh9sfXRPOgFWhHzMvGQNxQzDh
rgpcEb5heIJ/akS0En/oKYVioE+s19801XizaRwnmeUmrG6dpPVuTG8K6FxTS8Jv/c6oqG5lghR9
hirqu0WMtcp5/2oWYmEBOLAU2wr/SlCpo7l+0oj7FNbINxx/C8ue/K4kZEHtQxuDl80d5Lahsn4b
Fvh/sjUY3AJbJVzGaKG/i7CDdufALMfKq/k1qCA4owe6/Vi0oXJjiCnZWQS86mWiSe+wGNJ6/i9C
gFeCoyXszor+KvbRO9vyb7YCwODRTAxB+cO/zX/VpSIU3MjrzvaSM7A71Ubqj5q/pWjyJcB5JNLO
JXP42u0yanJCf+6LO++2ko1N45o8/lu6WUvlmtKl8tkxAcYDl8X+yA6x3yzkMV42DUoB2ZAhGtlw
yrFTFvCnaVtk1HBay+UHOjmDJA06djwoJ+yUSjA6Oyna6d7pCrjEBVFnZ9lI9GN/wtEn8Wpy8DsQ
Lt527VY5ZiFZjtSbxNL3DWSyUikI/xDqC//tKqd2NzFwrGyimfNydHD2h8n+yyFaehQ8ANeuadGL
f9OSiF85IV70gOTt+4jAy5zOYDZ8I6SzaerGiJaE+SzKgUuZPx6TrzmlbZlEKl3qILKSz+hLi5hd
Op5OYOzDYFhwAEZysP+nMe2gAlq+DSPJBX7NsHv2B6oaG+L55JvAQQ6+OgiYPxJwOVd9rXF/TTvK
h2lbfXLC9RR3/yca6KHrgIEIkIgJb1q4ECZZRwMKHLL+ZXaQQ8T2B3LU8xB8yDJ1+2FCZENO8HgV
lWHKoY41tIp4Z5zgV0PPwU6iEOyIHvEA7jVB/D1c5sjZGze0EEdHZ1oZ/tlzTzVpO2eCVnZzo0vy
6Zz2ajKv1SUy5vJ9KK6kv0k0DMRoRqcjOQwXLwOvxdsEP9Ww5uLvYUHGNL4X8j5YsqIE7qH8jzoe
ACb6hbozV7q4+NwqUao4J1FtOgy12Lpm3ps6JwwI9lARNFCB2gt6SlwSZVkSfQgLf+Kh1Dpdb/gl
yQvGTKZc1mM9mcCpHtab1i7V5raqCyN9XduKJKqdNwzWn2uicls9UBUeYHWsZ0HxOCEYTxeFYlaq
kXvhEpz8GSv8TwWE75uLajV3txSx4gAj9LAfqgH6Zj2VRhrzPMB+0PgwBSlL9oQkOtsVEQn06w37
BjCnIAs8IopNRgmfQTgSjbKrH38IbCp7DVDKlgK2gwkhGq5wmvvV+jbr4zUI5QlSJXWPO/bxr0Cn
wBNm3mLPMnhtche652hMMrZfIUOdLhRWLf9p+3sdeitHxBTh3FnO3PUP1QEishv4oS1SOjdFZwTz
1nAzdsQMqIA77pYPJscUImyhDSQYsD2iLO44SoH4H228Z8l4aoNqHl3HruqGDoN6LPHz/FyeH/j2
MuZHqebGNoHb6rrDlQiInnSxn5ZHWSlJKRpKqHlXcwp7yECG4X7BSOl05cW3J5hZlrZgtpOkXM8o
XHiEOrwxbPWwOSvqR8R90x04GIi4qVjna3891s5ssNRdAuKrk3smUkSbpkNeq8YOxmCq5v4VXU3A
7T+YP8VAZGFikoK2I1AaOQy+EZAd9tcPh4hZoRqMmfmkeke34xFNWYkrL2blvqwVM4+ws0gxXVUc
5CQdvomrzTZYXwa382108GFuJJeoTNr5d6He77xcjlur8F73zo+lX4c7NF4WlVyYLE31QCrPVS7q
/+xH2lO6QhRNBFU9BBZvGjMLvUEvh4fgxZ5XPbh0wdYuiPvhcTZ4ZRvb9COw/ADJ6u9Rs3ekiJ1F
KYMa3EsdqoS4L/UhVao2O1tv7YDs/WLDubzAvhvOFq2MV+qxk6nYPfajj9tvJJzeh/BWADorh/ji
PNsnwjWlb3xSwUJ1xIDDvvuwUEdfSjtdiYD80ijtxSRDYUPwnPMULkmaUe+o64ogLW56WPM9K/dF
AdZDDTrwHVJlf5jSJPTeZc6z43kuW9Y7fQuTVjZ55L0TAsVsqHuGkGrKGMO5/YWlG6Z4QEJHIlLg
xclXxPN1mkbVYfiZJBE4eOXLcWbCRo4muyHhtuBome1Nx0fX3MDCGHQAwMz/16WFhxcM97QOO2/d
6+4YhDLpMhmDjXpG8Op3rjw0uGsp+O9rJF3zp9q7DUmesV7YHfj2MXhXWQYMnCk1hOK3PMWb+UIx
NluSvBlNAlTlMzU370vBM6vUpKkhR/jidE2vosKU4EBLN+le5B9WvoI5TthVsu/y45OZsQDD/+Gz
hBX2WjBIAvYqwqgkf8Zls7pk58+/qh5h6Z1mqsCGW7lSikqAbNixDBW/zcYD2m92VYlG0bNpniFp
dOWLbGxqc5A7/CeliUESsKkg6UPnfJU+ryufcBgJW5jnpk6nFCX/cn6gBGNpRYpZwqgwhDacmqVu
m9JDZZ4shD3FWEvLS6r56W7t8bo16+NrtCOcvr2In1jMeRbgSWsrWTF3JjRZb+CT2DHmtyjpzzLs
E+agGRgzSaW3pbI8eZG1bKzkRETxduqHqIcZQLSADlPDaPxQ3JzV5hdw+OKHaplYVxeOa7eAYGdP
wEdrh6AiQ49Xqo5sjGmn1zImoUhTI77cm88WGMGoHS3lbor/a6U9nqNkGJJKJytIyx+EesbNItFX
2CHeZOQTYt4/s/9GEn7VA77FyF6rh4VJdQsEbqYxqXX9V29ff/A+9qjduV+QO0seZWI1IgOON8Tl
+mS0Bdat8lmJAS2JvDREkVT1OJre1k6f1zEz9CX+Bnj+eC/oYeSt/vYJ0TyECU6nKiEpEXvPUnQb
XfW1634ONskBWAvuVvE6gYF42FH/58mSzIVzrvfVELI6HLP/XLG0DpfED5aTlbmrVL5tEvJ7fSB+
+q8mGPq8cGBxWwU9+TR04dZ/HkooJTCF30aa8coJhcVoLf0XoWpsq0NYNlCmQhzZJYyNsQU64iE6
LG4RVV+7TsviUfOnp3xla0Ox+ZIbZVTzSf9VI+dqJcTamKBGq7eRxwYhroeg4W+rgwHrDou7gRkT
AgVKG/GqaukY4Lm2/vviyhgMLK7Yx9+Py+4iaFVjNtNZQDDs0X3dTN1GxwDpmQtXC3QVPVEKturC
6Ew8iehB06FqIlCHx83L1pIIcAQnmAgEk0+stPXLhOwGOi1uU319XWL8dY+kDchBn4VJHnK2dGCq
+FBrsKyslFV0rt22LEKHSCyTTIUMfaRKAGmxybByHWhmpIr/qjL6wrppwUgB2MYLaM1z3nnBBolV
jYQzle3HOwqJVWJsglyfCVQqFGBRgTxnqGsgVmAcc2cI42XoWIfJCGMG+u1RAXiHUPaMUx+bR+6k
9Q/AWnYhe0i4tXIyQTmy0yKRIaxGWbzwoATLAguavFv67p743xBirElxETUyq3a+Priw4Kf69nZw
qcv4m1FnkmWyiWv/9rnMal/NkFiTgmRD9/H6WtM6nTPVjlN4UBu3zvbQdlM5NEsWBfBBKw6yqJhP
927DjGXvDkOdNBmo/5BOTy7Zg8JgEvFxCmML/7JbA5X8MTv76oVW0NnlW04XEA/TIsHBoM5jGooO
t+okjIs9XpEzAUZ4yxrOwzNuCTc/a9JAxK+O79hNS4b7igvDo6rYoUaQO96NYwPaZO5TIVMSMqpB
MuNZp11X+BJyc0p+Kdp6MYLu0Fa3LxxVJ/k7oTTPBDYKFOM+usQBaBx0p7NT5Q+ZCQUkMTbTHBVz
nWISVcu9bEjR9nSCEEKz4gjUbIEbxI2i4t8nD2DPKVbvF2y3UheRxyl4Hw39j+wD/4O3AdP4ReO6
c2uMmbDiiABGBLF4JqNA5Xj2r4SlFGSOeAdYXKfkRiMN94+Tiktn6MLVVEwQFl1ZSJ3jPKu06eTZ
oyt7gl26p/qWvTZHo6BQ2EUPCUrZWfNxxb5Ws5AI9Bq1TGSnh1x8xDRI8Dl4x0xotxeHRuq0mwMm
9RUH/vEjgHSqPTkef3U0CqUODSn1KK6FUbnXkFx2vy4YfxzF0xeGMBKDwEaziHYylxLPuXKCmooQ
+3Y6x8eO0I5Go2BdAh0a46YtqJTH4U35kMRLgsZJByt+U5Lh1rTto7Yg5/8zaA6bm92IcG0421u9
P0soEBdBoxbtmj67fI1Muab5wuHodfi3ETGufczoDY54B356cUUDTJ7RX4qNIPZv9QDM060D6B9p
XxvMvTejiqNLxifh+/iQYPcq3b1nQ2wt3FTE/wxtLs5/irTlP1CunMxK8vWsUIrgYaJS4IAC90Cl
xs8hxMfSllHFIil4yqGCrvLjvTMCNf57cSIu4UGYbkOQVxQ6CVhOjUTc8yAJP3xtodyOd0Esqkgt
0tEp78+IJhDIvHGRUgvzmIjnEtKKdjtZg/jaGqDE3SOyYjsAdV8V0DtZSXJ+bUWHUcdcxcJadr3c
EE1W81aptFFw5anqaOMwqEn0R3c8NFL+dbo4fGfZuOr3Agyyfm1ahmD6MriAgC4R1fV5765InBAW
qgcxE4H06vB43ysFFnwGPL2rrv+QS03r8O/36ltT3ZWBD5sNPIdC3paEyv6rR9b0TV9uTtmTkl3Y
Nlb4eCgqO7aL/QWF7t40b0o86L16ziDJy8psnxyS1b7UecprHReUI42qhO5IQAfJ6QXeUHhuTRUL
Pj1KjtamHj4rUToeZGWPsM28KY/jTa3scJBxejlvcg5yAVMvH8CWizwf2dqFB/oRFtx0e8rhDCGn
c4G3Z7PZO2w/EsVv70rND690LB8jSnY6BMTUvIq3ArFuiUcJgGseUSduCgbfUTF2FFANlTiaZce6
jXQthUBgo/3GAgAWU6jta4gVH+xCiGEBUD1Y9o2gthr4n8vrkAGU9ndROsbCIpeKb4qNakCJiW9y
jZ2G/i2GAdNuS1MqOIv5+OVpcg1IzJIA5e6vY5sr0caho9/6aFeDsBpFOgCX5GRN9gTWQw0M9+fh
MwFw6MVGWtXY9yNva5CNhT0ZKRkiIgAkqCqzmSrZXBGwfh6mJs4Uhk2NSv/FDs7Pq2IQB43bdoqA
QP4ibZ61egRU6DcgW52WH4X2ncqPLeT61+REPSozk1HJnbdeBia8cEAqtIIOPOjC9i92M4p2sQzV
zix7BRVrTcP7zrrqINm8RmBpajHDkwDDuhWm6EXDSLJGT86y88fMrh+ANBm2TMu8Wuquq68obt+T
W5mG/SLxqofqH7Qcd1nZrcL/JkT4lvQr8Fe0xtQCowLn43F76bcAkTsmpva81mqIpkswc8kCt8zG
lbMDV1gCKuzO1WAMB058mnyDruoj/pgX5eF+OzBFz4iiIF11eZhYQq/geBjYwetpEh9K6PEYc2hm
ID0A8BaMLZ0naiuHymUnlAjOLXxiSodIudRkES0gY6jYqfa0s6glQSNMknzPIWs3NIS+aMbLyOZL
2RvnIB7lbf1npyMiuB7Pn3BTnEQdj7eWVOFSMb0SUuE8Mlbrwdu8yGUihOtQlyDhDktr15zGvxGT
vdzY2ORDo76vZl2PodpulIV8a7F8aaI6ts+y4CFMeIt3773FVaG4a+0/gQTyvjT6oH4jlUwFJzVI
LSyMhjMNkodobX6OY38qV4QzglerzAtkQgJh51gd6zXb6nlca0SPeJjxryW+HcyKEdoz+KP2X1VO
hieFZ99ygSX1t694idBWyyO0IH6itOP6pVbNOnoAU3He18mQ4QYUOksp3e5+XBH1TXMJjE/qE8ga
UvoMftduWhTlDpt+Q62VD7zP5hyZbQfJsQSt4gXgGzNx1uKFYU/QDZDLiDlmfCppB7micOWQDNVt
TJPBkAXO5w3EVX/3+v2C58Kk9aPc/BBTcmG+I0JDFcpwZrn1qv0dyiZ+ok84RO5qu6kdJPtZSjcV
ZyGrpUJulRycJans7JPkCLLzxDThSq+UeqaUN0xwrddxU4Dxs+B03pJzm4nw/yEbecfS6RexItD7
nOpd8p969zVpWIRSx0DTFaoc1q27TgWQPJJaF5azcOqJHS4mnAZb6aHY8Wtxw2BTbHioOuQ/HQnK
QHGbh5VPnqAoMKkr/rCFldh/e7lwrtP6CAmz8Bgja0UF+1yku6U073z8JX26/GKYpeHNguh6gQKj
sLrBJwTI+OogRftA8lGO3elJ94Wqyg9SrVY0IKorHSObPVG/vhiM1bF4M7iwYwgQ4/8nXFp6rYGU
Y1TUomCpEg9oJ6lMjdgy/xqdRkN73Ra+NI21YLBDiAQcfjSZuphmlIXuuYzytWS72lFgyOfT3IAO
s1YS3jBM/cFdq9ijNGo2xQJsUJS4klybVoWpw66X2q3msTmTSou9geJX1bIHQo2jB6WDaTtI6eVo
u1I2Wsg8eonB+BQHOzK7ljdx/ssaiGvIDucNAlDVzKKvnOjmPGpsMvbx6lYCqfozStVbVVdl394W
wBbD/qJvmr+6AqDU6JOWBeVD/k0drncFNny/UzDWoexjzqHj2tgewLwwTibRo+8t2I2sbt3GXEkZ
aInM/ClnWJo9GSLfRyf0Z2R4SWtla4GAQeX8v5FgdcHzKBhV7B2aNGrgjSptz4EVktm4O4mb3Oe6
AJ0Qlh6m1/rmUx1Db+99LVlSX7agS4vUZXhO3Sv2mUkApqMQNm7ITl13yF1z6dEVWCLxSJV97quX
+8Bs8m0+HvWl6GGcLujR7/FKlfAKOgKfQw6VP8uj5Sv/PsQJhdVvIeRx/v1+euLcfnxErdf7/+9F
29g2ULjZAUkbnR16Fc/VXMvEXZSaLpejKjrv+6gAsvDm59qlf7xAhorP7GNkUOLdwxo1tPDOPB/B
BtFpBEQ2xer7k2IkdGzNWPL3POWL0/ASnx1kwfF/vs4g3DMqA/4QBPORGivVdCTSQ+PEtKIzn7JV
kK4/Hhcqa+z2arsoFumF4vczc3/Ao2Jqg+8667yXmv2wwpE5CH+B4HxFbOn5oEq9CL95W+64wAuQ
BECttRNlvExPC1Q03yt/7ByHy92ivg7LtVGfYw4J7d9IGUF/Q0KFJohMn9p5nskrVHeUv2Um4VZK
rB5ciCBkkNaAlWLQXCoZqQi6SUqI28L43O/0W6utjHbbO+xYHnAYUdDUFyuwdCtjMPIM/tGD7wLA
ALTKK2nOp4IThx4W2+Q2wX5063t+eja7vCNtzRM7phGPSqujbo9GuS1UDsEezJniIQR2kQeA6dnj
dkuXMwUfX7SaBHYv1dh8kIuyM+2K0wWjyWmnROUT9+8mVxbHC+3vt/cJMfXmT/Gm6KViZ5wrnFZk
Lm1Glx4yFct9g0gJbhVicAEKYKGvtkwTBlpwna+nCI9F3Sbq65+ivzC25uwi3nLDdXG8JHA6ImdC
Lrc3VFSAlMng7wRSZzE1boYjWrYt+mE3rO93eN6lGf95fcmKfPtCG6fGQTyDdXr0rGq5Ep2c6WGp
RQ+OXzAuP8WSPpAQrr6Bp3v/f6ADMMM+ZrszbIdBLdUvSyCDGTQuRsHU2dYHaCEDH0aIcuy8/yn/
aC4m9tdLRGmeNmSex5sob+dytoXVUuPi3ec0lJ8U/Pw8MtHPkbkuKcbnpwCpSVhGCoS4PUjQG9yJ
Vv43ggrGs4R9HdKeJL1mVy7uju9K0rHt2UCsRIKREzOqU2L/XHFPmk57f5J+x132xbBdaGBYtS+5
tfMmFKtNI8aWQ7DfQYp/JqW5BE+V8CYrwUmC219dc/NB6fRbClcQN/YKQdq7AKKe4cJlxE2S9mAe
QOXvKqSaaAw5JI8y5L06ycaaaTnRhbGvUoxUZskWXFgF+Q3UHcrKb5lb5CQWp0HjbtDASOiYAZEJ
t+CxXf6tz5Ceb/ZgYv5vDn6DpMUV5HUVBgy4Ivc9QeOE8Al/AUiK1OEMDthtwuhZJhFayLBAWsBR
7FIGrBisguPKgekiRZMrJRa4fFTxpQkoFUyUsozsUamJfJdOdDbBChWdi/+2K3uqHXdnd1LxjQWl
wlJfWjbV7nnTatvcEZ0iTPXWkDGoDSY+xc1nu7Gcwtfkzx/PvQyv49eSQBMdE9mMWLNZd3CrjRNU
c9AparJuyrk0MszIMIZ1SWSf3Jq2+h7AaYH2h1VRZYAcPa/mmgdzEhJZw+4JvU+viR92rOvub4kV
xpC1H1fJDkLmH//iyvNoLJl3W5HSN6F/hfSuD435ZAr1/7YTMVYa2uBVVrc4F+LMF/+xD4EPWUuJ
uENta0hOe5N1L+3w/6NkBeGbskNm2YWhTq3IVCsGFFjA4AUAlvadeItwUubdlaNEp3DKy6CSdsLm
Ek55n2lYHwFG2MWlvAGorQl2kd1jmnSOLVmvYIBKxp5eTNc97l0JwQZ1OZpGZKlqZxeDMj9Rtzex
V/FKgC3/jt05zaHYHRWn83NpEj1Bq/F+uNWzQtBsn/glMR/8UM+stI3oWcx7KicKFIUvYYVjqkA/
6pr3szB4wRzMLPqTa9H59Y86gjiMl5cD1cFmpSPDxy77KtqbLdb0OILuBm3eMU46nOElp6PMYD4c
vzr/LVH+bzAG8ncvAPxzIWVBB8ppoZIuf90P+Tk15SCEn7gl9IHMH6g9Ng9uAStOdvvOiH2S4X8G
ch5buR812Sa2clat3K/aR2ikV3tPWuggxiVDaAFFbwrTTfQf84ILTibuj3PAWyy657USKdx79RBd
KSkQsNCCN7mqehTS6Cxp0EkFMD5v/NgQt+NQn3LacXB0/ISjVYoIcVGNz1FzewHKDdKyaOpU237n
x5Pxk7HX/v+reCfMgq0d7VVdTuFiKKzbGVFop7kDMrdBaeAmMTLx7f/vb/Ky5s2hg+/HzOvj0tph
Z1hN65rFjh48q+uPmbPpcH/vqrClXz+lAEDSDnIbb/sH4WRXzmFKSQKU5gqCzNHH29YG6ZlCifiq
hfWN9whVTAD6m4ZwOo0B33p7ReIuX53WsbdiSDGlGPah3Bt6c3xokM4E07yxj9FQZEXvUHifTRST
I/kX49VM8wktF6d2F7Icw5ptKkoY3wukqtLd/Ehoih2k7qCOxSIDwWgy/WUxisNHJBI/M4xLoURV
RIYDwi8iR9v2DdI4dNSrAFEX4SORa5Eaf7UCy69NfFp8Kx3ixccbvSd+UucWM6yq9l1Mj3SwJl5w
k2z9kX5W3zl7Ik2w+WCwQ075m6qr/cbOemh/t+HIX/vCKm/Duz3EH+83UcOsjeB6Z2HvWZ3minFU
lIa/Dkh2qKqhv83l1+yBkkNMwjZaYGZJMj/lVWDupRXg0V6vcEFioxr5UI6MccjzpWddNnZiQpP8
bvmMmcmmw/6GnZFHPyqlr4qK8iOG51mdIxmgg7lwxSwbZEwHZUiOaXn9dEKfZzZplBT2mrAqOvVI
bSO94KkmYdb48KTZCgCA7WyypJdS0lvhiHsQ9SFeThPHNGtsnqzgR1tWVuicdA0++IA+zySE1h/V
8Zom5AV8nU53KAurydvAWnPGLUirKzr/UxrTfbQ5mFpW+W8aO3+pd4Io5ABgmZKOh2IUE6FOSg7X
hoLpSupRDQw1t9vxeAYZcEXrPIbyF2GutDoFWBVB/c83xyDLBHk6eSGKiEOr7pwc77AjWl48UHbL
xMg84dSH23xB5ausAM5L66GShV2iMKSa+EQlt3QHkKRf93YBURO91plphxxHSZNq9wqbO0Gixg4D
yYeniPamOi6cMnNfl3pgU80JDeRJObjOfHz5qXc4UV7dD8kMkZp13jLH+732/8TmJMSdVMr0BPHe
6nUi8KnO1UbvjM2/V9CF1bB4qsZh0SUK0HASLTVo27M7y1MedxI6NvjI1+QQsIja6KBBQ95RqPx0
bcaCUMSrad157Jg0QUquXQpimbf4Mx2K2aPZhYwfud02RN3XpcZBKvgV4kLjDp/5AU0nPqFkL44Y
ddTwOvuN2qjswIaJqJEbL2Yxlmo1ekDTSLgvgD3HI8QySQCv85akA62/dug43r2C6FdMdpHTNEu+
Pd3E76ovIqB4BKiN9ul8j/mlyMw0F2ouTC7irv4kIESx89ivbZzSkhGlGJNCC6MUtxT2wAvzV+4i
h24Ogo2s1cymxSGdRbUYZ+OmpWfYzIfykDa9/lpo1uPZdUYdLVhaHKedw8Rt9zFUhp6+C3JQljnk
VXHuKAa1pS00q+rLKwUSLxcrEEXUUGiYZULLJgw/WH1EjQVt8X1743XRFRk+PDh2YpEauop7bG9p
9HYY5y0ZXdPtnfFbivs7EC5F0Nl7Cy7N5kgfzpPxa8+i4rBQfsdJj19deRBxug+oi1EQhOVamLiC
PIXqXjo75iqNokGuYEla4cLZPo4P0e7xO3M7alDjdpR8FVrWjs3I0l28EDYQhWcvLSllyRb5lOuQ
pJdsy8EaSbVBmvzZ4gMXj2+HRcG/mtD0gGeHAEsV751svXWI374/yu1wrzOifGSVIbB1Kvc7BYd6
5LpGh+TQERKg/60rM7G/TRbppc5nlqtQRwrYllCKBxyYkhGfISpo5avUIFmUdsFLWJh2EZrqzoLJ
9f4kV7Op8TXqLWBeardHmgr8BOy8GK/jzhn9OkTTOqlLyiZXN2N9CkUEmqLgLTOIBrNkavuIuKG0
aww/Luf9C/OIUkNP6VIxNwikMfCBF9zaqfXrk2QUcJpMFUN06kO2VBLfkF6khqYfYX2ZnCYybgCJ
46wMlQBYEGdfeAFmucdRmLimThNyqU+AUIj2mRHMnDrUxUl6p5g2ngWcrze4cfj4y1plFUdLL7wt
7Zmrhq3BcHecfqzfbE+dtCP26nM/uKktY7PWgx7i326i/oJgQiWYqrGaHsFzQ9buxRTYdPB36Bzh
aeSreKS7W7eBkqH3sbQ8YdgRcnVqmquhTkWuhTgqceH+NknKpwAu9iiNW0QgSZk4eE3qpc6krusK
9n7a8sAzuPM1F4BVJEKYjLvmuriRrKOJ0/ADJhg4G9Tarsc/7IUdMpbqk0tvRVYAE2kzp75eOw9Y
R68VuLW0dHU5kPWzaGfO5dPDRDh8qV83OlN/fU+8LbMHPhBcBTDrEnVgTg6RuyXcXVInNztRc2Ni
opvF8yUSFnTga+jXtN7a/HSG4NFzaqenmhlBiFREfEoqYRwoRbXXgcR+RtdoKcQ8iagvJGH2i29/
uyTfinzveq5Bumh1XGZ17uoN+gYGbv8mYHJE/R35q4iZg5pGpVLoV7sMjbSzBJAJuhaP/U7GEfxJ
PMq21qrvFi3+GDqoo/Rdyf5CdepRx1eZRd13oJtMXsrnT0nGqz92p/Jxo0WTkr4zd/4XcyGgtfQZ
XIdgLOYCezuk+dsur4MW75D7DDPhh0gSahGtG+Ux/ZKyMNub6CxvNSRlkNDLpqfl25rm/3op0WVq
RJbP1ak+5OzNTQkRA44Lxrd8/Ibm3KEv67EP/+5Nk4Be3xhM4qOzBkAfLAFjV1pQrBGufAV9uEDJ
rx4eFgujzhzFKE2+vq3tFs0UK34/gt4uQJNyCfGJXsDFsR/nF9GndSJiWgmUt6TF9zWljiCH8c11
mYSGiqtVJduhe3OqIv+5iSVxDvSQt1a4BGiX+dEUTgrMlWQEBwHEly8/0MIH/qUIaPfEn1br1CYU
e4F0l3Th4UPeIbagcBMVZ5W1dNM0nezUB34N1VR1A2gM2471OgxUw549jOvyoy4E38x/+1fvkv0a
SwAputZlO1/1O4SlQCLrg1iGreJ+zUYBasbV71FOTmZrASHd5y+rtOtpaEgi5Q9ft0ACR9yR5dXu
yPa3v9MW32Cp0o6qUnz/QkLSSl97uHQYW37Wq7X8467BHlyUH+jQKspGkVT5nQxPfvane/+KJkj8
yxMDvk7ONMblWLTlabnlHju4INw10FPR2d0JI+hyzfLJm2M5s0t/53sUMQcrj17Au2SLdkYta3nZ
2QvYnPSaSoV/xaUPWCY8Gv0AOxkU8Uc3oCtGTp06Qo1L96BwqtZwBkcO5wRJqf5r4MB1q9JPM6bR
GmhV+a7+LPltT3JY34mUcHXKX8iZdZ/s6FWqcxZ/2x2FHlawP7EE00OiYtR2tyiia/EgipIYZYN9
qOBh2JkXn7uZNHYb/RGE8M8BMZa/Dfq32bYXnkg4XpctqyM8aG9KnHHGPKQ/+fuDydqFPFAyBKwL
zDTU/2C8A8laDAMGl0392r3illoe7ZOxpelb+nkZNPNTxcx3Yvv+JtXgMhbuKSK7/iIZ+eXQBVGs
maAnOzwCFRaGRnhgr+37xK1VUh+ypa+sEen67ZA7mvXDipqCTlklQgVht9Oh4ZtnNJ1mlCFgQiV8
v1ml+oPbWzN/ZmWEcUjnx7JC7VkdZN44H/18b1ZxAIX51wqF1GhKX8ynFKJdSctT6eaIHzO3wlMq
4963pu5Q/Sdt+hULDuBrZFj87R6JbPG7G2aTGebAdjphj94P5N1b2tJ66ARPz5Ta/BUCuMDbd/9Q
1IopSGc4m+5gW7YYcYs0LSNcVOlTnScYimWQjaVGSCyA0IhCtDnM74Z6o38M5fX0DCd9C6KIrtP8
eCT2WaNHKuZy/TcEtuI7WCuGdRUx8O3XHBwzYKEfCdC8AqN7EauGFA19QigwNqUjcMDTYvxZQkwu
SFmUeMSlB/ZDvlNse0i7lA3qWZ9KvARLdotILpxYQe4/9nLW7DwzrYA9Tk+jtjprq7FcC9TTqqcH
o8lo91tFBEjIJAfEnwHUTZSGs9dUUEJOY0v6OgBMvNsdifAOrhQuANHl1sCnG0+fe/42WTPyfzhY
hpiMtr5j5j5kuH3nYnt3JzrLCkrgkTBot1aS6wi1ugEG3hjt6vGq1w7oYTHw9asGCsC4DZw+EXPD
HNUQKKgFb2SRSKAN9fdnXnfmNg89uizTfvBrzf22KiOLI3oTQnH0pil8gNpNsgF/cWPIteTTuzTC
4e4I/xJy2moPWbM5hxcFuPcOqvgSOr/lkyGkosv2ZrGuMsnYZj19nbTgqGibhIwyuDCZv0bB5PEx
qfoqDAjm6aMhUA9VFtrjodPZ2UI/FUYBPLJ7yfl40QmRp1TxtyUhGSmhq4KR9CmEfh2RgcQKZGK0
gBtywa5KKB9yszo5PuDKKe1RmoPQrD91wTpEjnTuCsCDMBM27y7mdrpQsrslSuUYVwwyn3b7VDJr
ZKFTyfjTlG88caAZvM0/pfiWABpiS+BKADGQC8qRwgO/itU6lw57dT8W3s96rgww+bbpLl2MQSb8
ECy4PuUU9HgCIhOyjUmDdMjWK2diZF8pfEUhrKnpkhmojUDPdFfXdloolcOcNa1EPstC1TJsQcFq
cfRDFFxKx9fbhak88T6Z+RQI+NsMBQIZmWGz2q17zx1zq0698hzHv0OKQtWF5F3SE5bRbBoqM71W
yAU9j9I3sVforicpqe/RPmBNmxKm8HD5ce3WxaGItg2keEEbe2PE4vxuCe84Xsas6txFTEUdrJdQ
vdnrlqh3F5yXAgtz/O3VcWCYLaSEC9hD7qfSHMLQAU1SrYjo7gdFLgRPjFIy69rFTmpgpJ5Trwqf
w27a9xBXP5ECUj5bFyLiPS2g8ms1LsSHfnD82bDwJKU/ZxCCyWOXDKSOgvIUY5MyPxSHKvUfH4I/
q0xPKSkNtXREYu+h1AACZrIsvJ4ACaXsTaUmEjUxMLH7H8fbc0Lvt+RItqv34OabhTeQa4skXkbQ
Jdj2+uWBGmo0i0WfrkVlJZBjyx8Ix/8ySJwTybcwPBvauXJGqdmX2CvEFzXIc6fGY9VdvDiu5OSA
Xk6ZloZqijsuT+Fns1pNWRIR/L2Cag5bzIv/9KxXXO6av5EXFBZOd+LoQwT3P7PHng/IFtXcaVvF
jWSZEOUjz/spGv7FsJO77QbJOhOnOuJwm4pkGBidtI3FfHFdDMfjzIwF6wVScjFaRZus3JFZEN3b
8K/WBUO4rifLPDWuNC9RUh4TAOYRBz1rGEK3YNp8KkejnwoXei2WyQOWZNR7+Ftl5ecOpO9eLVAY
94vIkCHLWsGwwq99P1EoXiGE49M1H6HEowoODvNLnxzes5EJjoU877Ig5jUOK5H+mOnd+OSRUdMe
gP1k7J4qOXRXlz1gD8WEAwbFlJSVsSFllaubQP5A9ifOs2DEzXCFqNsluSGN7vmqrQqwvwO/9gjH
ch8qMV7ziWl3sF3lW4w0z/YZMETiup09IVECXvrHoW9lHXG6JcMrmy2/2SEJgdWp/mhLdhvf2Ib/
lIATMxDBL+MViPhgVp0t+HLchgHqQlo4HR/A20qCdHn3eKYSPjwRfz+B1DcWJ/yH0W74uP7F9nXP
DlZZSgSR68WwPK3Njvk9NHU7t8cfCIj0Sj3CZOLdIVimdQB94eyCuocgSxB+ndLHZu6NLhAXzDuP
qaoD+fUEj7B1btzUI763jUmgc9d675/kudLVCfUSAeu7FluV76Sz9+x1IIIZczXQ/tVt7Jnoxv8o
WGaYYTWu+DOEVf60hXT/t0g8J1JVBcfXWvyVVClXF9+hobNYaylWj7xDKhLhn0YsLt22m20Gw1OM
owErViiRDMMZhGFm6LGeeWOTFbbvXGslFz4lhM87wX963oPFyUVbIqiPPzqvaClN6yFWLoN2qFdH
HJp0VyGFTldS1VtZLVjd3NXOwy3Zb9CTi9a8WjgyUYk1ZmBPl/xtWTlq+JaSAufjx6yWNWS2j9Uj
pxOe8PrYtfdWnEsn1G2bjwC5jAOl6pRsKTLVImOCk8M9OiQyh7CbDslhXsTOKRS+Ra2pC0KBa5x+
Kn6VCgreYbxuvXZO/0+BWcJefwBwd9wMmZetgXlgH1zJrgiA8l5VRU1K0XHwhnkvPWg2bWNjFeIS
rmALaUyA3PrYahvYr0c8RbvwZLit6/XH+gIKc56uxO1KXYiAPiVbLndnPkxmtxtJVO0ODve6LNEI
ncEbZ/g1ozzQnDhu4MUQjFgQBRyJsOsxn/lrf1HQh6ghmpPIxIeTMR6RHVeil0gSN8Ddo7YR1Vbe
vPYufKgr1pciG5lNrx7mFmjF6M/umiSo4tosXNdYnJkmVk5BhEmqMAmvjaE+o9UgtD9j+Ri3CkOS
evoT9aiCBCF1+o6aW1RZ1BErgWOcKUY8pYBlc3o3QcRpKdWFRLaEDqTvH86zLHyQ5ntnznRGu97H
DJFsvVdxEBF8BSmgJ9BYnEuJdBukhIvMlLbtqfGGDYsQA4N8hJXVDK7yD9kni+d7yvbbDRGeMafy
zaQhaphGFBszZyuPQEjX2deJ6JioVep4ylki2R08tXRmTbBt+ZHeq4fFddRDxXBJBjBvhhXNuRNB
luybkaKVS2mfXpDF1yil+lOOVVH23MtCxqgV7NBgadXcHVmYZymTN7qZOK57W1ima2iVBcRTFo3J
1oUesU8DBeNveQLaZwnrLXhVJjWEWGgoMgRwNH7GbX9R8Xk29ka5nwkeOTN3lC1ni76qvqIzRlAD
PD3zANuBcmRbWl3kkij8VYqKH6ULVYc/tuzR0Zh0cCtMH9lucgdFwLEkYKSDC78F/GieBScuDdcS
meX/3i3T3lDZ897o8Nxvxwc6g9ybet7kkkfBhHJ3gqRMEBVGhwVFCJjZYkUsUlqvj9H6neO+3vDr
rESk+gRoyHAonzZhxi8EzCn/ywzl6TMd6JzNp5x3HhAI0MiYN+z77wtV8tDrLAlszZmd5/doboYk
4sixjRAcT5wcS3smE14vTXUFIFvdv2YbpQIeb/eyhaOPlAgpeGVm4gaNfRsaQScYfHB5Jc0odYo3
duztWaTkvmcPu3ce1ZS07NsUMZ52QhNWy5uq6DQTZagXe1WvE8+/z1s4sz++iPG8qyYfFReevVq1
I7TpSsKxjm3QeZqhBpLABc0rKCiLOLfX/eQmLRPpHT8LIUidUOWez+XMGMYeu576UmjbICqLYbvy
7ea9SGROwNnw4oRfvw6b0rTMOVfLomxjujRg+6rQwYsqbo1Nc6drInDEO/YLdzu1K2t7JSAOhhPE
8NG40Yo1jtJwKGOh60QgqO4E+kqVDuxtqBYGR0zUHyn+yKJ+95s4r715d4KblChdnYYGmv+DxZrE
z6+ajUiW/vKYMj6MMh+3/rQNMxn4ptiaOPW1dKh9EHwArbcpsU2vVk4A99RVUSp2b5cTdB5sz4im
g+wcm821R8Oiqwck7UtuWD6wjT14/3gVaeAeiOSVTqVg5yCHTWzCefczP2lsjhSgZl4A/x+gOuBu
1+DvobfPdtTG0GwEzBq+pgtasEqOL5DDTOW43ZUkhnyXsD7MTEqss+fyKkApVxSDHuq2B7+uYUrJ
alpsLSq2n4pvjVtlAR3oSIfYtSuDdzyyif2nxpeqjA/ColsEE/l1vsIue7jDVUKuG3L3V0ISNn5F
IKQ0xuJm9YvuW6vN+u86QlyZ6xFbX6/zSWSS+iDvlTgxVdU9HWVD1wlDr4F1BMFUYE+QCO/htVrU
J6mt3/i8MHDAyyizMHvdSDGghmww0pIZtzp3d8ScSSOocKISP+NffDHpSSikZ3WJ/0BkqgQ+C2OX
4SseuQNaaf3GPfLsG3AJvNwf25zTb/QVaHPLGusxfILo76KW75VXmPmYV6FPg6XEcLx0qkB5+NGu
Z1DQYx4PiVwgGXPqfACyakfVRHj4AtxfeRzIwMTYPmWdjjBfpWLDsrtRvWLHT9y+lRZUun/nhLox
j5RMrzHrlg9Z5xvdVUWMUSMVbYwMZ0B6hprT7Olxwq0qds1OkoEZKVfvTVbVDqAKGECQn1oWNlSn
cUnBHThAyk0BpYFuk4I4hoa4c3cdoXGhYYtWHy744+R9afkVK7MD/bVMiP4gdtqqQDF875ey2/pD
YdNDA+ClYwZbJdVgDRFkJgnbDw3+++xim4b79kbMubuu96zT8qgH88TU1uLkXhWTjnN8Wl2X2roj
m9EOC5B0l9xq7vUTGQWGGp3j4HpimXIXEglraXBkE+bHIk3Q5xAe+vEoqTqNB7vpftR9LaYBD/uY
COE21F+xTxByVtT29KK81F2qgXFwq+Zv0c6xzJoIHmq9AcexRouZ8AiPnxsHbRk3+v40ttdntPtc
A+VfRFXNVh8uIisEh2HqDDPHG2iyoM5vqB+9Oyh0ThVHJX67iV9RhUxnu7mxPSvw6rvAMxUFN4Zj
67LWG7c/RQdK+MHghr/p19GSHT7gIP0dy91wY6OKX92OHury8uanP03O9tihxe/0epCeAAbL4T3K
2iLRyi4RNP/V2qJbDAGK35BkKXY9S54N9tDgDgpsT9xZsd8J64oHhu8wvTusT7R3Pqh6CMy6YHO6
xUHur7YoL/TvwIMtXe7RtU7S+s7+lr9XWuYY+vXCDIYYEH6kaKAXOZQbO+Xi2ddYBRo5aaXVVJG3
R3FWgb4zJ8mfp3QNHVdkduWACgN4zY00eXXZp0uTe70BfM8iCh3eQ8PKoAMgI2L81LBvrcLtZWpG
hZlEp/u5NAA08VY4Akx2LM8+jO16Yu4yMU22itt/My9A2pc0zINSAT2uSLYMI10WtVF52hEBzBH4
H5p10QT/+WTzPMy+PqmF5M+1YueCMT4BL8Ej+uqUvq7YWFdigOtz1E7demJbm8jUexl6B2DHlSA4
c2CkBBTR5Ox+MldAgLfdkXYKm0/65ApNA7M4qrJsDUg8EU2dBZxRUVhdL2+Nwnh9mrULtTLvW8F1
Q1XOaYBZvzBhOL9A7T7W3P7YyNnf6mZL+85vxV9QT+3+ZUoN+xtqsSZEdAyGkOyd4XnEDe//kQZZ
KDcq/TUKtaXWzoPinnJcNzNZhQmNKklYenwQeh3bNbrihPqGfdd2mfTNem2iwOyZvAWwqHFnRN81
j7PlI9ITLZB0EczSoJAISzpt/XaJOPId8D4AVnxjbAzvoS9JT1ny3LDoHlWHVGQ3ULgjPBpEm0s/
z+io2xsXKyEgQCE/zR79nGAQM2vbS8IQdLYrkaJIc2RmwcKtulYF5nvws+jIYzQYwdJ15/pv/YRf
MXAqOvYvlw05ecTwL1hu27Ez44Wht7Yad+oFz4yfM9KNrkI/Cg5HslhqszUvpa8wjQ4MHnxRNFNs
p+UPUc+chqt+4uexZ/QA+PSWkafKvQewqzZP+J5Vef5+5lMQVPqY6Qjn+5gpoqX3P2EOOW/OkBFF
3zwF4D5Pwqla0QMk/aP08R0jZf0uDuKStxljHPuT8s48fz3b+0TPuUg2UGXRAzcReYMoyVqB1lYP
03qqVMQTEZ90Rj4t5OW+edF4IzO0oNJnMwvklRC0eXRr4n049fbqrL3W6MfySMQxajPvlPvw5Uou
HgV/9qiQsSAkFtrU9FCytXsCSRJitNpTqDTTq4deqw71xhZlz89ho9UyqK1u9+mAZrRrAsIk0JJ2
36qV1IU5HX+NaozkHLZwJi+drr9gg0YE5fdUPxIqaJBbz9jryHjOq/HyvmWp2SVnVeLfaBSQoLOs
k+2zdMDOHMZcZmfobPZc8fFTNsE6Yruj2BiuJZd19WyUBcim8NvHfNYr59UUfb5VMn2wlesYoE0Z
rq8v1XUBTrKk8MN3fiBs5rhygZG2bG8jt2FguhS/lyQkRhByQecVrwNEQMhyIvEvan+nI7pTVqNm
0alRBtFyZQh9fXd4aJxtQvIO3Z8tXwKWbp3j8MX/6wtzjmdi2LZo+TqFv0JUp3fhPW5nUZCI8rJ1
dZdRyjZwo/YF7cPXJm0QiZrPzMq8W2AvEO5/3B+b1DtfYpm34z2B0xDsQ/J28UYYVsChj+SOdLuH
GtGfE6jynResW/MkG7Q1ee/rG8adojk8xJR2ioV0yiasK4toAYbz4cpFqqy2zdJn5Wiop5mzJz3W
jfpqtYSYy6+3IL2eVRkiljNwWmF8aEWLIj4WbRQg604sCLonGCG/2RqSgrCQnv8cP/233FWqQgTb
AdenZRVRuNApb6Gt4RPwCKti9p1Lr9J4e8WhgtZfJq4i5aqsUJlC+y2q0VrpKFV8eRibxd0vTnY6
dGq24rd0RIRp+lWEELO+HYmf4mSwKJg0ZGJgNNLM2Hsj3ko3VgEs1l1BomIrTs1VAnQSrOw9GaY4
yFhcoltP09CIdGbww468JQ95vRZbGFKXQc5cVcLn2VSWknX+lweHdK8SxQzqrBA/zAGUD+3sBZUW
HVsuK0qzAJ8F7Sn1vkZBuwysZC0PXtTxzAElarmu3rDhH47IDWtbfECf+LUU1EUjSZNQf+AdXhci
7O5JAoHLIGphkyPVBXXbxFyFWORJ3DCtumuimyj0pntofJmSeOJvRjxY/LvK2lAo1SK5TJm+3UJf
G/6xP+kxOv4buQRC2JgXBOq7lsoi8RYe8Ews54Oo4Trb4Xrme2EJsk2Y3WyqmETIz7qaAeWRuLe3
cjOFGCLAhaq+GAYTmYUnkfnccUZSGcWzhTCr9LUyh5EFcYNX001ERMqC4ar8ECTyuW7hC63HacfB
9S2SfgbqmN+mlPYHwE7Otb+35hyS/Id3o7q2XHPMOs6KxPFhhonZMwy7DoSOBTW+alrC6jTnXT+m
1YN6JI9aFLA1aaAGJC+oXKL24Uk2G6YmlJX+THHu8QqsBC3m1BX4VYmwShk9LjeFzIfU+ncmpqOO
pvzeAcVufa446l1D+7pfO8iDjt6hjNhreFMwN8rajGgubOb9I9SpYZEl0/eHkzDpRYJvXzQOdR1v
r9HmvgoNI+bpl4tH3vrlQc+NFiAKl1psPLWns9hOXbXwURU5YXEx1ourfKrAoTOqyPshjjvasy4V
s2WYIYRZYqZ3L/Sw68aVlRu1+qvHN066OKI6o+PehgBVvhSIbLs+8XAOK5FFLBlnUamzLsOUobCC
CX8mcNDU9JYEAWEaamTsr/Z2aseekXkZUJwRMY5nwh/+lLNFXtc86aIpqzgOe7rHeGmX/BE0ure5
LR3WQN6b81/SdNIVyVmIezpHlCknJFpYgG2rtgWBNnCRPVfyvC/OmQCj9Gow2GnTuUN/AWa2CF80
IYb2ettfSbLf2Fgh69Bnioy+QQkWR0tAByAojlLleTL2w1JrDwa4Tya+yx32OHOH7h71x6B8elmC
kc8gbFpG5tboPFfhER2sCmYeiKFIPGXbR+yezaxoCfCP3nG2weZIqPYRLNqnBhLuHra3AkVJ163j
NMUUNtbsQ6yv7mgqp/kTUghk18Culo56Ssb5uqf1fOIy+T866zvoCgLWoFiGSnfhDvCTLj1b8mOc
3LhcbLot7A6CSciD7IFyhHzx8aVgboVmMYEklaj6UIPDd91h1RBt4wWdYNN7W49Wt90QYJwfJtqp
NNErJ+WndRC1ZFR1eyZ7okwzVLrCM0VDEh6qJIxLeY+xltJKv7exW1TwP4WeYwiJZNjyXhO6jotQ
1ZHlSK0iJ/64c1xWdfPyM4wnaSb9cwPqxbzuHcljqMc71GEqDmf3WcGLHENSOZDgZ4+QsUqqEvKI
/OaWrNkIb88TiW/FJC3OIFJjyOKBiUp+Rs1KVfblaMDFEViZLYO/Z278W0tHRklqYMk60B1iuPuc
e4GZ1Gl95d+guu61WA1gFyb/sz26mEq71BBhG9Vcz2f6/durkuXBoQOHMr/NhQR+32j7MK2NeGTG
r8sgUW4IR/8oGqpOd8vYJMp0IQ1Nu9brODGUfvJzIrVkkM1vI9oDNmRMlvBNww6xy+7gzdc3PqP+
pbYtElNaIjhcZS0UlzoQAUTPqmfGbQslYhd+9U5wkkpPFgzJSqKpl0E8XAd3A1/jlC0oipOwXkiH
5XlbqZxNE9groXCzuDgArr7RcmZueO7V1TelFEsjwrzm3kc01kSUtYpzJ+c+OBp0xqfkybKy4dao
nAh62W/z7l6p9dWAdDbXYP7MB6MumHmiPHTlJ8pY1XnJg2RwmuqYXMqJTekYrkyS7yTQU1a28x3B
0EvxSHGF06GrQCZRkCv+cdUF+sbgOzVKFPQLia9e5SkFjV/ny+rsTUND16sLPifQxZ51Cwogszyu
XBJUILJrJSkn2ez3ShzqICax5hbIvhlFFbblt3xWicwRyClejWnSRQWn/Ps5HJ9++c5nmu1Fp1Jh
DZanLvud5HWdsU1TwoK122gjZH+Gr3MhBgcL6YJtR48LQ/iprCb8ftnEOubRL8VKDtpwBbI7QkCx
wPBWkeb5wePDlBoMcCPYOstSSqtHOzrLCL3TXihVYXjncMnrF/OujTQ1y736bJc84Hp1rzmh0U1n
bQGjonW8ogA7SW4hX3S76Qs8dmWFVfQQ/7Z0afFr00WiFNEh13OjNnYV4l4Wsu1Mz+oc2sBiEqU1
MVmtXQoyU3+umTX00eYOEPzeZmXDZavfABvJjQICfqOXzMmA3vm5DubU5SdxC8mdwZ8iN31TJ30B
s9u7YWsnUbANK8qupUS6Q99mOE+R+ZSL9MgE5HhLj7GkF2G/gbFIB7zAVRRmXwfbJen+nHZDELoH
7GO1bnUulraplEP4n0ALuRa+ZJVDQjoE31V93kepja4rkVppM52wdiDZaQMziMyxWXq/2laL7i/k
MjlAXkWXcstAcPEiRETVCE0plo7fTmsbYZ1Go61OyNetbngpWVpT/wrPMzyiUgQm/yF4rqi4o6UH
jSQSlbw7+kYtf8c0Mzy/+8bSmgVbWezUOfU6EkQM2SRiJCxjQIOKy0nEWmwdpnblAwyJvFnjzf9f
v5yEYSQ0u0aLOUKj5q2f7Zm8qcd05Uihlf6+G1het0gKPgGwFoGC35vGl5oyfrrKWJGW4XVcQY4m
RDZMG5ElGoASOGLVfa66aMAH3CU2tv7sBw43vpRLpHJ+xKElVz+mcGojTEsCLpkalUw2+k7zezGC
YKA4w3fqQX3KjuSoF6E93kEXgw5UKm7z92c4W58ifCRCy5KlundEaITir6F7lpmYXCjuBdqsY54n
XWBDnjB4iCtGvlVSRwbhlvTSEAln8Ywy5scLRcQJP7RFgPG4Z8QQt9Jpt8a40h12M3TdP389FZ9a
w3NcEDQrwxUB7i9QiQ0WPn8RicULU/C2XwV6JtOswywWfzoNkqa/vLaouh9l0oy3ZVK/md6/6D9z
phPTWpo6MQ28/UpPkl/a9NmQvY2n6D6UrWhhVGHQ1dGltWVr8idQVtrvXH6pRUEjS3NONygyXTsD
tJmrM4tzn6kK+gpq5HCIuYrVTPcSmEz5yaN5isxyYpse+29GvOSrFNEIQKX/5Y6YIxRqVOSLS7Nj
0AT4nEuSBsldkQyRH6eA4oSGv9K2mtJ3k1NzVtRhEa9k+LKkrqSDBLGjdWUVGVtnVh1CQmE+KbYU
4NnNxx22bWhAuulhFcW+nVuN+rfseku1yCFnrhWeVoneb4r2WYih51XsQSAVJqyS3S9gU1unRS91
faGjNHrgduq9hEIFAVhuLU5u6zuZjSIxQCnHCINOdRGx61l7FFxAq0TFUWAT4OMehrhC4I5taKaI
nABd56IrNIR0QxXM0OolWRioVIsCeV7XtwlaDdJBcu1rSEa9YYSDnssjDv3BEg63qG6oNLGPXO0H
nR6xDsskx/3Frx4w/RIoupq8qcBVkEH7BHRoHgbbGI2Bwgm9kHQ1D6Kmoby+8jW6BCewSwsZx0dG
h8eeZxBwQVDItduSkAIumb4P/oZuB3+EjQa69h2vn+i1K9RWRn+BXE8JnpKczdP59fgtGD6Rpivj
j4Vx9mfgh6ow03jOVVlAKmjrHTzQgBcjbY7PzvxH/H3k3AgAeT4xFyukpo8V31KIHp+t5ppj2+yF
YFoJniUtUS7fcQKt2vtj3XSfZQqz9D5IcAL/Tn/NnKY17EZ06KNrngBU1+LrEj+ItBNXIGuTWFyD
T/reBSYCqg41vhP2+dXwiP5dvujG2ornB9iLp9HJMGYJOX9L/Ip+MB0GnfPISPwflO/yEmfpk1/v
omnGMqTLjWfHZSlrz3MKedQjTTsSf+xbbeqABcQ2sQCPqGjNYNZgjiODCX8G3mkOPL9WvqjV6Rbi
Zldoxgsm0aXcmWaxSm7w1QyZDnIE5n0nCVgkE2W6wKJmpi/K1ZcPlkRJfXWeH3EcyhzWNamHpKjV
rpw1nZ5BFddR7bhZG/ci6Vf/lqMF5cASbyo7ArUijo4RWE/KWAYERqp6msPwBDMmQfO4RWX51zDi
4hC0iHYrW9MLgm6lV9Xx0vImp8K+F+9hmtPhBnVQQYYU2V/afuzzf2IsL4gm3KjXon2ZLP343g4Q
zSVixV5NI/iV/a/JEZRzFpLlFK7UupNSQDLm5Q6PK1CIxwCUpoGdLlQHEKu2t7nnNjvzz8nN3BtR
aOqgx6lyhu7XqsfJkzHNpTl8LVvs9BWmsi9Zsnamyo0fqz/l/QNCz9z4KQrzX8y7dspGltBpHzhk
rLBzoOVv+8t9FoSA0HY7U4a+q/nH/IXAJRhTsPthRLcUcDmqA9DiCtG6/wXCmzjIXnoutogOMhmP
74y3kx6GCZeS639kHU8MrdJvx2cJuS2lJ0S3aOMEnBtaIFH06NTKrY8erioyVv7vJE/meTBjfE3G
D9H5JZtxJeu6FURw+sDQPp4bgFaq6paTG014opx3CRiqoHbYV/rWAD6Zb5AmQpjPkfzeoGdAtu/x
xM+6Lg9oOdJ/0CAo50TQxddAmN1Ki3WyglIHzNOYUv1GucaVFxXsy0wewFglreDftvwy+Ql5EZ05
wcNSnAgiv6bbCOoJdPgIigyKKGg1CMrhpG+TBQBTx8vrYJDWNqdyj1+O0xIXxGLiorhrT3ZpPx0Z
eQjCI2VB7uTJvAWXh5k8NuTycscqNRF1W/50gkPtg6lhBH2OO/sjzmGoBMhL0ZN5SEyqzpk+zVHs
NNNBdloZfOJinrHuRAqsSlBYJcqB0p0oODGcKMY6CVlBWMPo3wOsqkUnyC5l915EI0t+jIHZA6IZ
XLggveEQlGs6DawWA08jZ3xLj3gehzr4XFh2//lGbUnhoMU+syvtU/626yvuXi+x90Cec4pXFc7Z
zk1gxGKp7mON9EehsU2PxLpPbzziq8OXf8qbuGP/HzcXu30OaA7w/lqylw7Fg2z0IHt4ggKkPBOP
QA5ZFXJx9LvtlTZACIQZUabeX4WzjnEvDGFOd4u5MMENxADsRQNSgCBPA1edPHicnbmgA0UGcMLg
15ag8iU1Qjz3VanTaYLbuF7mIgodJ663UbLHuPsBLBRayg0AUEf5DQVcjKWd8utsNfbPZzgf3AAs
P2KEu4iJTBGIqah/UM8KoA1fl32pUa0I/MzHTLArdK/gzVmPxZR5inGqZFig0exiDkSCVs96/XXL
Al36WBAttRVCHmgXqHknbXe6jOiGPfdMgRD3HIgRWv+LLDcS9OGgFAfnTE63DpZ8DWhf9YWNAbHk
8fk/pwyLGUMIYk1ognr8PVpRuADZYz7DYPkJP3wXAeRtrhpmzMvo9jILwZ0SDLzUW/2ij873lx1H
Htjw4EftqTIQHpM5jTSR8u7CmGyV/SLc2JIoixmGPm22ayQU4pS795LWhDZv6M/TOJJlnpi9VB/I
S03JvNuGcENuPCwddXyKzVNcCU1QvAtVjCvht75LKTXitrY8l0ipLVffuuvSuXaWUxfweXNWOK+j
StocD410iILQVceTUWn1tNkQtYuR+XARVMKyYBZh/DWa8ohIEctRy/4PoTUvRi62cSS447bpDNpa
iBSVEgApsdzkaVrIMtqwUvCo5qhOV+6E4zIIDU5ZEJhJfqjkTBz0146E/y9yizqGc/9UlPl45yz1
p/dtSgU/LkqBZnjXpOlFytMOGImfaVMDblpYootlsoYlnlHdyPX0yrKmxMgG5QZd59IjWG9wfDlb
L9TdPNnVaWPesB+tE6vQxz1QyherDLVRyrzB/9a+wsX448Qoy0zlApeEaQIfUTq6WQOkQHGeKS0S
ih7sT4Mwro0AFBrqzjYWJl7cuzDdfBXGmviQyAP5+syJ15HabMfCDxhakDIW3FEwbRwwIcwfoUEe
ebmaqfPC0NHwkTYvxMV1aX4a5GArQb23K5Wg/4fElUwWEDmYeXHiaapQPEWQA9mHGx/djIl6J//+
kq4GG0YqShvEV61KPax7hw6CZlTpUpgPI1/xeqUF3sYhMsW3+Yy/n74gooBH6uGRUVOeHy3LkDT7
45+jQ4cvZlc3sR3JnlbMLjJxLEUEz5mGgNO5AxUc8XgOptx63pyLA5d/HmdraS4dspe7TO5YH6oO
RSfSuMFxntUY10kTHAFdFC0Ay3RJRlJ5IC6FF1drcHfxDCYYsD+5Sfo8ccvYhzbjlkZpeDmvFTH0
Obr95Ca29LimPuG4Hg6NIZO4gdRR2OrO/pIbu8XVUAEl7AT3YfPHQaciVjOGa+wfSSVaGE7255mj
9CGFRrhyEa/iV69qhufwISesBLbCwTO6ZrlxAm5HbbYm3nL4qXoLGETL1q0RHfP9PCwt8kV4FkxV
DjggBqOjnHzZKHMvQuNG/IdKztat3p1XBsoAYRYIkvXbKkUo/qzTkUnruablRkXxuBD59x3W61eG
qLkUp9/zUsDJU3cjJ1QTC77IBtgtlVbSKnq2dgciWODMmxo3kwu5Eq9YgvzxlihqO6u9r8m5Q0I/
h2AFKDRY6EgVEW7ejPu0UKxQSATaWpOoBUFt6B1LRBa0KN0pmnz6Hpr+Ly3BSV9ZqPlbS89btVL2
kyPbZMNDpSx03081DvHLudsbWK+VhX6YzgVjY5dC+r5KrnHHf45YyVKoxRyzI/mDuE0q65X9XqxR
Y4hau4BR6y0lXXMUVxslM6kPXnAIEGvgmu6uYDA9/yZYyrEAesDrk8bYVhcOZbInUfqIfx2w5e3p
fCP6RXmiBTTTLtFX+/gYc2kpkCSOg4XW0Nqfj/Uswco2Fcx946SR3fUEJYcJnpo1Ph8Wvb6PEk+j
2r12CemEuOEU2JgAwlFqgU+cOtyRQR9NRTrlqpONLHOKHGnn3gqggLoSU/pm87ZOV+jfFe7sxhwU
ZNgsaUBGHt1OiJj8PO8Qb8NIUVhjomAJZBX+f17WzPFHAN2yEy0W6cCLK/yd1jnu+5+SThrAlk6G
30mRVaPUN9AG0PnUQ0QDApQ7mEekqgy8HTd0yJJyX2A91I+3xMXt6Adh/ZkqPMSNCKxXWbuPjJyx
e3fFC2j5AEMjs1bbDLLlWBt0GvHBXI6YqEJbto46U8Y22254qCQM4D98niYOeqmXYqsJ91+BOTm7
izQ5k2MnA2c8F2TLZzPTLr6AnkJdPjeeq1p7gtTe8RvdYGO9t+TghBPBmUpQ2aplaQOdJhw1gnQk
oGA1loN90muEcSqgmRFHzFbBDL1ATujMAb0Hsj9/dxxl5xHCRhZktO9HifuPpO6Iqre7Dtg6pwOu
zngcO6itEeBWYBdu8BwdonLP7oGdab2LKAoayQ9LOnKH5EKUySH7z5LwYQEFdYUzXVSJ9FCoBb5V
qTSO9moK0dMlh0niDup+9x6d5BOqk+TxFAso0wDsgj7ATbZLaZhNwO10T3Seflyza+q97FOe8EG2
PmCX9LVcTTfaLG0IOTqqB4HsCI+wgSOTRuB5BwvN+RWXrbQccJetweEpV0bACWZV0DBHq4nMgjfP
aRHxvhotzyC7Osmt+RoO7svBShG2BhXy88tvvViSVCWq31pfGanoc2PsOVxRZ8D6TKP5GdWdJvaz
6NwHeUqscDBO+6l8ua/z7f51VlI+tZiR0CudqkZvmbN92xzuOHP8H4jhg8va7g0/RryWyDlQNMLM
1lwEOPIewQ8A7AvpOJ0RFXOpxOoMJHY+cOe0udZNNdsDU4z5wCaf1I2nAlbWMUY8rLzl0CTjZar6
lT7WjEC+lIYLvpskyNSIbqrRb31mn8qrRt8S1gVKvH4SHDQrckzTM6vOCS+TpweslaMukLM3wFMb
6NHjZhlv5AG5pRs64oIb7fPE2WjTtJEDbEK+nEpj39vOk7osucChz4iuVRaKN+2TXSlD2qQ8BOOl
Y0TxgbColbrjxTDbg0yOOEq+xUskSZM2tdmZhSWHIfXP8+TEDp5t80DzkSO0BssGeu0THVnuXMM3
j8p78Qu6J9gbXfeMLdUUqdmdxuPYcl1GuAfIA98d5vQhe3K17OVC5H1f7RhbdbD6IKP6XwdR3tBJ
Mc/3yC/1UsqoQO9dId1QgBBYiCC4osYeXwFF2ee51U1wUShz6gjeUdtuUHOAhSGtp0AhcgANzQj2
uh4STT7NWbqcpwArpq23jGpkDuJbBybHEfAm1vzaShIVj3IOcE8WCW/ncZ3MkD3cXl3skhT6aZ9g
lnDF1dZcj+D063beex627MLxHr010bSfo+m9sayg4V4uQrCUyMlnFbEP6EWiVMJaa+LawHhjXJa7
Dk58DaPeXOywZnxGJA5oygfy2IZJBMa5sT7aGkvVK2hOZ5JeBth+q8Ex491LK6pKiJZ2nE2NTUs5
h5jLr1IhEqTuFzfmShbxcCyA96ozWREnEWLwbfWQX5edpj35ATgqTJ+38/GlcvDLtOWK/n3HiQlk
yyqaGcx2hY4aQwQ8XE3P209ppLopnG9ca+k6Yo9UGuX76Wvph+E6g92xfN2ze369+ZIQ0bHQIKU+
2ahMh+DQFvH0onbKn81k9JRCAlwT9+v4G+PdDAGpYQOKPvJCTw9t6ts6VebL001fBcBGV9K2APHL
iTHeOXCS6hDRVLZIn8m56nfsmTFqgETDqGd9UPgRqrzgHnhJmNAwqn7wFiaF7Gbj/WVOHFr5tErO
ockfSmaTVVj6q6H2SYYzNWZ9b1zCHWHRp0tX9aDDU+HB4TgfTqzBVMy+fBuRSoop5DWY17Yfp8P6
X164q6TNI6Egjp9ik/Q/yeLfA4cTkJXzxeRs/iviNAwrBIJPaxluU65uppK4qLc0HX+6OeR5UR2f
k1jzRRHlZwZidMGcZkFle3mhQM/7pRrl9d9DREIKh0x4K+gFcEVYUVwjas5nLWgYAtmX1QIIxcSt
afm/2yCzIQnFlfwk6vp/LlXnsl37CLdZMDwCI6YzKlZ2jyxeMdVXBZDclCItZ9gkne1jcWAA//e2
b6t9PuHEBImUAmveuddevwjfmJ+rQldW0fUcR+aCp2jIskmOLNprGpbgrp+RCBnHeOz6owYfT1bA
xjlGS4cnxH7OQhv53rouTclQzq6628PT7m5umfKZcOwoBdROLIRqHXv5Xu968ZNlCXw3XybWaJlK
r3/1GImZ7G/kknwnEIIykrD8LekZiS/iGauUb7sdUzuYrCqwB7QrSoq8+YSj79HmbXucVpuCu+KI
z5dfLw9juqxWR0QQDt99cAOXPoRBCMPck6dBs36JAH35kL/IfvLn74sB7rgScdhRuF/59A5eKpeK
vHrX1jlMkyw+3rIni7oZYllNpAvHj7lwumSJ8BLnDi+Yg7y4HPKzYnZC1BUBhlxe7Fz3AlXXiYzo
5QxLfHKeh4uKin3AZ8Vh6J+BN4hZ1Q9WrbAmJ2hbVxe8RZdgC0LGRM3KgiVJNym9ox+PNYQjAGSY
01oulREsbHRxph0oaj9FXxTsSo7GelHrnikqpMGtukpHhVCDj/FvN2BAbrC1UWPZOT9yTc3ErUfd
47bOG5omGUUgubcSWm9TOtfRDHmCInHxVtgBBEQyxbSTera/M2SeeKTBNi+4zYx073fJTYpEgDlu
TPxkjYPeqp74EUQepE8v3w9waNOGXUqFjmK70FNOEieemfMI13OepzBOCQHwUwIJmEkWSMNgT0bs
bruret88mh2lpdrmU2xERPep7dGCyFL2yWfM28nUQylZ+wyT0Li8UjfYirv6oZT7iqg/P+XUs7En
w24XJYpPq4IFao/EzpflkEfnDiWuMBWyH3etkbCRZ6DlpVqEMpWYP+G8ElLPoGX2P9/EUo+Kfkz9
iDna5cOrqx3e6ZWzijFl/NdbbokaUyyqfQxPZiGuXjnd+RXL2fB81lsyWL+o7pYeqlT9P91yJgLr
YP6WqCMLgo/yOpS6U2KGhmYrwbq4UH/+MLjOX+AiVITtUIIJxSmlkrj+Jpivhb/Ny16yz3xPpcgb
oWlMib5S6qyPz/BEVRQAE5P2f9DaaJl4iQpIcjqg6tMJG8DJn3QJI4zFST4jU+sXxcrMJiRla0h5
VdCxfsQULY9OhUCOwgH+6P1/2l/Ka+N0+fjetModbiPIFq3bZj3Y4kqhaX84FA/EAI+L1uNXo2lv
ocatYgrtZa37bx//dn20Fshbu2i1XKoP2vQGyIuDMahCCOmZJPGFjq81qdurjFoDZaACHPdz2vlC
efIdanswUdyn0eJyDvUXCRJW1ObHKnljkAIX9H3Uvi9XW/rkyGBxX4KSXQvKiUj43JpXMHhKmkSb
UeJu6SDZe0dGFsP6afwEEPpcxOCny3wHIJj+3J9TIWIg4TX9KG4r2/oZWejRYr3N8AqPkSgs3ic2
HqWi54q7k8KBqm7idWDhEJpN2IcCJtZgZYDg1pvYe4Ew1/HEzpyRTEt9K0IcS+hPTUQsVTm6IE9h
mlTcSeSNF825wdTH/oEGdsVti3+mGNeZsEJ8e8YlIXvuYu4UpqcR/0sX8XNOM1A8X6EeE7XCAWfS
hkOn3JgTMqa/3ouUeEDbEdGeYWHnRvjFvmH9yk6yJrwQ717pz+s7mDpkJwA8RVvgRe5vfy15pmn7
tBre9kfJvGdUuu0Tn201DjWlKo0fcbbr3sJs6cMKByANSv6ONTiS6NoKBzpvgBwScpNZ3r7LqRAE
3hT728iBmt7ni/HTlnEqv5XW5QN/ANQWEnEbTll9OyxOMBMrfoDUKts7cfYthdQIosR6r7Sh18w5
E+RCNOMkC9FpkXSQyHaZBrl5ZZ9XWMpEKvjA+taTaSGe5Po3QnFj29G9ouFv5ND+MmWhmCg8nmyK
79KdfO5J5KgGfIo8+2xGFX7yCBzx7FFZMltO00lJ/idMRKU7Owp8Lezd8K09/PZ0GEG/S8nnOwdA
dsnB+wGOYJMjpDcfzd6Ou5yCGNQ/1I3OyuFRqCdUA2+S8FsvWAMbxcvN1nP4Hz7yLYb0yICMoG6I
YHYGkMDqOql9hHSxwqGnJ+7LRyhudlw3zq46u+DOglSdzlWGtJxku/8AjewgNw18icx8A8ImoVhG
c73CXnNf8DwiwX85jjjBIvE7QXv4IvBmGX7uo1GB9P9c3ifpkgKEvdQ91xth2pAo0LgdpBMjxSqE
q+xRsQIjxJTwte+A4W+A9mpwOcdtFZEX9InhzmHiIIX7iVcrOpfV2aZU+NyviyqeEZRBVPN4Acp6
xganEG+XC1z5ka9Vw/vSg1uWtdw0uyBTcoqSAj78mymNbN9nfo0sQ7NLnUmfv+CfyQMD0LOdZWwv
5BwHD7rWVZb4C4DSpck0Z1YRih4kEr6apib/rW5CdnE8vugHXGu/KtmxNF2zdptVrGOeAhg4ZXH/
k1A0Qi0Rg9CoX9MhbN1ANvRGTzQKOM+Tb1a8hbNPkCYUyB3zTGzeIGuvuj/JZGSxftWH/ZAtCCjg
Gj8JwGK5OPThwiWcR16gp62HOdbj6BLSL7KWvRPlldnnQy3d5bMDwE5nrnQzgWBHp4MM5TuOh7rG
fQRk32df2HHhoR+Gm6lVofMX0wyKdVfhQK4i3VQX1WY5YswirHlHV0zJOuTKwSPDp346yj9enqjz
j/wZpTqYyigL30Ic7iCWX5NqhCxzt8xGr/2cV4tZutE5Zw/aBg64JdABd4Uq06aDnZN8negIpTMe
WkNLEGWZ3ElvS6lm7igj2fvm/xo9ECUf4D16MQHXv/lm+tmZ5jzT1eQJuWfz3Wo2gEVywojb4dnC
+x8fCsIhgvm9WzOejhsHKlHHwU2PI7YTjP9BVxkH24+WcvW4Erfi8DL9G1zGiFdjcjbA3N1vt/22
7egAKqhfr9tA3qsfkoaO43c0T/kC+lyZdXHIdPa5vYlGlsDJKHdV77l8jyYy3iLIlURx05Ks0iz9
bXDpYERukc5gz2J2PWoMomTzCwaOVeq9XYczwkEvd3HtMCy7ZBOp6mK32ryqrLuyqE3jyUsgqIxe
+u/JrvBc3zLe6vUklb8SMKog9HQ3IiyDwjNlN05yi69iRFwFs4aGOyxFube7wfkZLQZC6qWh+QxM
m+kaCfI/+FZZlAdmZoNh45uVIbZS87HCcj8byysLJsHB1KCnOsXWKvlrYeqC1A2uoVKkcQsOF591
453l5nUnf0ejR+523iuZxjhH8r2zTQ7wzL+mVnJYnOjTpaTPl7QenOSWMeCMtQn8wXgPBqmp3aqG
HV8CVwAPe0R/u255C4TqvIDUskJl9k1jf99q8vIOKZQPu8vfC8JEHmQm/Wxr1+4BR07QaqFTwlAL
NEXEsAO9UD8GAds9gBf9VZkXCvLPLge+CvmlfTfcF0hogr4zhIWSqzlPhhrFifoRz16VTVd/ceSI
qBQddkiOMvl+QITXLtq7In7nPfbTVVVEJ+k0HErFUypNwoIHiHtzPrEhrBz9mSIWN+FDyNajGJLp
8/pjUnH5ikDCAmb7NK5OfesNz4d9oSOsl+tHH4jHA3xa5qyj/Q9mLHn3pc285TBO2tRqL7LGt28R
wqXBLCb61TqGKQLm/wRBnkdbASrtWuNwDZQUt40N3oBFYrfYwCP6WNfpO8v8j6mXvru6gwZ3A8Ee
lkNvPKeNcH57fghZiaL5Nq+beIM3uvcRYoBp1WXznEZgfEEZ/LktVlUoK7dkuP16vO51oEq9+vSw
nsinLTQEiuGtSQKB+0vQHFcIXO69B5FDmPAAQRRdxzxWMThWTMBiCDJUbdmkcE32dNkKt2ehzDJO
AaakhZghNn83CQGY1Q5qtHUwzP6C8D83HSu2FcvuooGQKC8eZ4VXCIYnQxbQqsRBNP+wyJQMeqIa
1ioUQyo2gAtc4fC/tx2w2X/pHa3AZ7adE4IPP81QprvapQI7bQZ6T/zOcPVkMbTRELqbAVDDCfqX
j6wntOxtKCJLYin3fbHg8LaBEq/JJyPxBYjurn1YcoCMw8yyPgKQ+Uc4MdsJT69VVg+WPOYsXY9s
BjZ+Hs2S7Q1v/UX3ehOsQL1vJNthJucRG79sSXhqS0o5msuZK2880rBUB7S3k+BlTHyMgnlEMlRF
Y4hun9UFl0v0QfBlairCxNmVpiymh8zEXoHfdMOubTKONJdvnis5R1GP0PxJXPZYanAYkCIkKgx5
p6Qpbeuj7jbfmL0g7dJEd1e3zA1fHbvFoT3wMSDuL7yd0ShCaT1S+gS+PfBt4OYfNy5yvEFT6nuP
8Brmt/dxQ0IioDEBUrbzIm1ey5FCs3iIe5UrqSZ9xkYZljaGQjgq2KNU2xNCIm7HSbPdnoIidCo8
VIc1AOTK3J9In52CK7ZNfj4W1EzdSLdaqMfapIlkXfmP0o8IyO6y6SjublN7A19o7UqtWKugWHXf
KlAVY/x2G29WwQpZGB6jpjSLLqIe/kHBOlh10WHQMJC31TbFwcyMLR/5Ehi0IPuABdyk+4ZPrZad
gJSHtqs/DvgiBOSB0wk5IXjEilPRhbXNRAdNvWMlBq7xP2tT7zhjxBsWyIJIlDzwDJpY8pigVe4k
kkB5fwAO00sHGI/apxpvzrp96YdDC8ABE0/vlSqs9gaJ4hRC3OF60JQLec6rwWBZvV+X5HJx5VIp
Vv+Nt05WXWp2VMv2ydRp03RzjMW++PYxOo/1IX0vwzFKRZoKkYUQ12Uc2tEwyMfzlp2/apozMIuX
uSmEMWprY7+YQMaRd3GxGQoIQxqi8MpMjkpVcvMow5t1Ck7yqsozWH85cDgSRgv5iNGKmiVW3/5K
oXMNW+0f/o5nC5qT7hCGP30AzufBhtcOucnvWcVUyC/EAuBAimncCJNIuUJqefwZZKLARoePwL+W
Dgaq5b1FL5v0O/kmUQeDTTSl+GHofE2buwl7hzYj9BK6eSTuA5kFhkIitPz/vk1mhGu2qGxscyZo
7yjxuLjDZY5PfhGUC1CL0epT9op6rDNkgXHjXPLvSFRKPUet6fKistjPrMkhqasUO8xAc32a5gbo
Y4lhFH5OvV+DW3KAcbTnv2qk9QiUibaFjJ0si4ubVSCX6sOHHNYL5N8tDdnNbNT4VNB1NH2ZYYEY
ds1zbABX7C/zpC0EadELjjo9uT51zWUIoZXiENDGC+DUzqK0YizKp3+GHVF0UtBrLsr06PpTs05z
O3b121ct+wvO22J9ZdOu59FpsqCKjMHxPLYCV2LhjJhAdwD55nles9QUpJLM4d4iH2a4MAhSGQCR
qMQcwmI2oX9qREwyHb59fZibMdEd4B592X+Y+ZrbrXX2rQzAnB5izXMLjHPXeDPw9xQtOB2hUYF8
HGt+T/TA95afHLsVelVdpNDIB6KfHHTOyHXUuUySK+rXDZMJOeDcFqgIVrS0WdP6N1w/Kaypl7yR
AabeB+Iy25lgzgsg2Wgm54CwVJ6uIhDUzD4zECtcWszs9Ykd3dBmD99xzaOKaEUoDxmUPWba8KIP
M3vtDtTxvQe35xec3tUw/qB5PEwRV7uFFOO8q+ttG6gS6wwSKgIjMNkZYeZtGKrz3WzjZwS05lgU
P1KCh4MT93SOgO+K7rTsBe4yzm31X6M3XjVQQWrCAVDIHRq/rLLv5lBMXhrMAcEsFlNEOCyzwEsG
wUcus4GGTENe/V/y0/1EW4regwGFg/srGZdWM88EZXAg1dcnxYDBudc/JuK0ZqdSwB8yw61bthQa
DZEK5fwHBBTPCus7Dx5LZHQTRMad46Kxt2Q2Uc+HB9etlpzRi7PzsGVZcvZ3Q+2hiQshdPAgDK/l
NO2+skan2eEs8aFRZxY2WiV1Dvcgw4+KknS7hw7yLBXQaLuuvOQdMxI72UE0LW3jsLyVH/kmKcwj
34YU8luvuZDa4hmLy/LAjJoKc1qSbPXf+VhQHTiEqR/QNetjNKF92zyYuAHirOMJQuq7GcZf1pFA
FUBcS/kmhmWifB0dUsZiUmKxZSVyxOqtn/7Fj5QPaJK9HOyVuMC5GDXZsdq1lpWzzq9usjW6zmsY
eV3/zAOqwebbYUk/nTQPbOQ3DH30yPBJK66TQjmJM1+CowLIYTcz2ayqB4jnfJXWSsOvDnDzxfJt
zN2OHmmwo9qYb7XJ/6XH07RuxrXUEfc8D3qKgcuEyGUQ1NXtvbMSgUkgRjiIkVEbDyjp7tGcWfFL
5UfWZCcJx7C62U6qz+QhXk9F/AsYXNoJw9AFEF+/OFKpEhuR6PetXSFQW0J23oQ2fK+Ky2ZxPA9b
dVmIwZCBm1Ga8VaRG8ZfgKxREAQVHvv1wH+0NhucEdkiE+GGTjSScGhuimBSPhZdEwaHUQYk0MtO
87LXRlKg6797+fLY0hgZ96xJQFTmdSd02Jv4YKLQlo5Om/mTTvMyA1uFGFERvo4Z3CyS2EozYW5m
YlLCrSRgrYFiGpIVYdyUUfwUf3G0e0N7Uqc0n2YJu2XUZOf5AOdTbN0LL5qpc4tQPBXsxhW1QGf0
nUpI7AUQeXgiM6JLCbTZzCOUEzegoSWgUtsJ5t1fRQobt28K61IkJWt92VA5NYz/N3uKW78QK1+B
F3mkI0eKhDLzJMfTj+Xt24tkrjqFJ76uUNo1hEQuLB0yoZk1Ja5GjryLs3NR+QnpHtQr6zfi3kbp
2gy7cfnES9YGo+KpMGZ+viXrSJGQ4/guL0M1W3P2ynutwr83Tl6UcvPbn5yXOz58lWr8lreHjQJy
DBkL9V6bn53z+SHLUkqhEYUnMUKeKn9q+IQMRytJeP9M19rwpQS77DjQZwc4l/XPRjZELnMTfbWR
68pX6Dy7Xqq/AiWjhykXSg9nB/2L2wvHVkjNYBJss2J3SRBlWZn1PV7Ppq7/BwQHiqwVk2iMO0V+
eo47NsPK2RkI+SdG6pcU+UK88aNs6TpsrC3gnbiskmuAFO1B3j/Fc3qpAviRVLgX8sC/PKXABZew
u5Pds3eYP6LcEnOJX/51X56nrZoL/+5Urncp/IR7PjELYDXGua2P1liXbi6QQf7f4bMP4mI7/uBG
3YDtbaQK7fwChQVSQGDtQeW2cx/Vep0D2VhIsZPdN/MKeODe/G3+pfPofX+LSyXe20RpuKVdOzR3
Ho14PWCqfRarr+1ebX5eI2Wx/45H5yoeZ7YYad/GwlLeLOUdUVojm+qAveRY9WhcsdLOmFLUil+s
mfIl3OyL8WXMXRiGY6bvzchQ+ToYpynx8bhElzzEAKCbKzOPaFyC/ci3KiPYGOSfy+YBn8JBZ/Au
bkqmxjE/GoppQYh/Rg44COd+LNAXHYXzX1bJCvMsivjeJXbZRRKEqXlDM9PtwbaZfHVzPKCLYy+a
oAGFgIZp46hub8+BLso1wkN9pErKUEvzxqkO2ahVQ68QWvKIUf3mCRzFCkSLFnneHB/Z5DZ2lS83
kIV6cTRcLgIzPHTWtHSYOpwaf3IgLdWxgScDtMhz7ZK/AV57pwxjeshzGpnLN83Ask0ud4e6lIgl
z5rpSVnvLpLaMaIr9u+XShda2wHLL3FUCCFpdZfks1eZ4BYvaYi0//25s5/HxoEns93Z4MNwQSoR
EDOCBWxlf9suiV4KrQHKSagi4K+gaf9FTZ05OpfKYqWW87VPJ+8NV++agTTeUvtQzhXBxFYp8NnR
fTZMgtpSxpun9e1IjaLtAs1fpEyT0aTTnJDNAVYvdisAwJ4weik1M42NiRpuR/SvNKTv+mbTq0f1
zvxwVyxgkj3OXMpJ/QdDW6mgF4zacvcObZy8Lcxbi7/91IanKTSSVDyVjk5iribCjwbzvXQd4WpH
5KgkD+lEfLjM+DPCdw2JnzckaQ73D7Wq19TcWm6eKz3PHj18DisxgiQnJ6e5S+/CCWrgret49opV
ufFp3Ri1JavLvxHRNRZmmE4Mr9VPEFtdg0RLR0jcrmP4YCP2Uu/sme8DNNKV1DSzryRpU+iAK5jS
16qZFXLEQJt+OQDvPJ/nCqc2gcOLfxOVmPs1wM0hm8b3e5FJ/iSVfIplg5WglGuYmK54QM3fx+Ig
9VYdymx481lQbyL33l6mJ1kBGs27OfkTay64puI8mNqd9FfOu/4m3AE44rfdB2iVsdfPmV/C+Biv
ya8ayJQsOHcpQq/rSHmkH6PRRM+kdrvOBLWPR7mKctH6G/iErU5FJX/nrtRj1CxoeqWAgSnLpsyl
Mqg3dJMvYRpkRe0XKsqP9M7uPN6qyo6sqSDJxPJPMos/+8fqCjv0jejtorVrd09GDVRxLpKd4dUx
SQuoKW03AouKrPgRpfUYcrVSNWJdPcpxzsNgJYbcBTrhp1D2cPQBcNCxptmhNOJt6+ydDEKy/pZZ
XAkVIHdJaGcDCFntygS0t5sF0ksqXmJy+pkrJVw50MTMao/V3U6IuWhswXomVqjmRSqHfN/TemlN
9Zp4ZFsQgcDaYMsj/BPbgqp5XzCS8xs0taB9BZcfViyQVCj5EHynY2QuGNedlJm5iEYG12yuWVc4
ylrK1hlDNxX4CerBtXQBYCqKRyiOJgiokOPvPXBu6v0gKgxFp36vK/yGqBGZpzNK/S9tF1cQmAMi
xrzQUaJklv/RxEB73OtIPM8lLTKD4s3kh7vGuCyH7sES7UIhXuZCMxQ8FG6drEXesiLjeFIpEeN7
xU4l29DOvg8AwrDtRqhGJB0pg9VGHW4fdCztNNljTnWcw00I3y8Pt/zwvtVRf0cLT9pMPhCvtEe/
AfdsC0WLPCGWNw8oAiWD0qgSUR8ooKAKt8lZseYqyXyj2YbnPHO95CBcRD/RMZsPj/WIiorX0+7Q
INeoB2f082iPtmPIHSehczNFd1Ezki676hXI2az2CTZQlcCC1bT1E4Dk/Y2tXsNIgEgMx1hGCK0B
Ha0jDkUdKX4QRC6fhkOtkrV7HlxsRfMKFbEwWXpwQfw5pXCvljoxSGJt/3ptKH/beOEe0tEe0WjT
FlKdzUIRbg3GZ/cd7+BVGXsyc9hE+prUvP+K4vfHEI3Eq+AbTtRrIl6R4gZ2OK9cHfR701aNSJMG
pQGbUgFu451fHF9e7WvkMDpTTSFm0xxuplZqjUMk4QNbKaVoLZw5uyJ92/WL+uw2R2wIilSLFPj6
ejt2aaw+LKFXuvW/SNgsrECufMmllAGrFSf0tmksyinSK02KkTAZudhbl3gdzoXj4HCSlj35bsWj
OHtGc3mulNr7S8T2dFo826XZkafYIx8lJgK5pnid6BxV3lHg2UCWY8K8LoUnvWLxAKZdIN2cV3Wb
rAnF0GUt5z7nOD9Un+EWBaxYdx/8FUQht8cLV5BYZXraWEy6EANlwnBxU0HVut4XAeXNFjQu5xNZ
+8b02ryh6rjIqSgt/uNwk4AWPm+hKeDGMaI78rJrYZwCDGrgvHaxdch+afzyCDR17mcP+RTH/5Yo
LGWGy4PijRFSK7QmoEN8oo8fHvLIf1vuwOuX8D+3yak05K5A9rBe2xgYz/VGBf4ec9FLoob7MAwC
DuD5oj7IlGhUYyDLPQD+nc/ebd3WXsoHiPxXPdk31MnWpRQxNGjMB2yEPM61h301e9ulx2loIxOR
unyQsqXz7n5fyftsB06sthVX2Kb1lqhsO7C0Bn2T5Lf7IfkFRQExHiuPk0/6OFEtKr2gKOZQpZYW
vuUQDUzNrn7Yfg/kZsoiqQViR/ctFocoqm+rG2YAEy/QfOtQwn8VYjw/fYTpLSulJ+Cjpy+WYh/d
mYSsTPU9g5K2CpyRTITKFwjuBcctt+qymU540gd5SsXQ5DLpj+OP2eM1m4//lIx9KS2+5vIJueps
OC/gV5dHEw2Qmy9t8bAszNISC05a9iRtKTuwt4ZVUOSbT4Q4PKzrHyZY2H4R3H7LxZimz6h0mwkq
EZPG+TDv34HtkaHSg8Q5gZ59/x2ecgi005t/dNmOEwo+jcNuMe8al2BvNyq0mb7qG9kiPOpwRWtO
e/Azxfy5kRto2A57rpu/7m2SjXKMgRzrDYCwtq98iSB6Yces1xad4mhnjaKq+7KnBwEbBVYruD6E
eG4a0q8X8jBoRBl29KaapCmzLnJ3d/dQA9yUt774h2bZhXC0zus4gS/m56pYlA9mcwBMKh9tdJzD
TVpacCLnA0F4CBWBJ6GInqf4kAn8k8tSrusCvEpN0S9WqI4MMtw2Vck7bdvs4PBffSWrSwhd7U5C
m5qPYb2xVeMJgOtheT0zhPaL+E38DvfgBpUgDxMi+Pn6DovTJwleaShN/tPIz49RBWrYCnlMAADs
zpjUY4EkAv1zRmAGNSgBEkWPx2OqGPSTPsXzwHKlgsOZJ8D+t+lF3tHT+bT5uoszD5aLtiGPE6Ye
9qMtMtu4y+IR6T+nPqGxG9w4D/b6cXJrcE4cUB2ipLNBqSh2Xx4oRJOzLSTpJosIJicJ3m3FBCn/
JbhF118ljWf6A08mylclM9Mvses34jwPWVZsNmlD4RxeRSXfjLRLziiuY0As3zVmJA62R3bYpoSY
x0B/gLm+Dq6kotqU8auyA11OKTbh1DzTKXeR4ohBVu71lG0NT4ivKEwmK86yft/5anxsqjH1o5xj
L1RSBEdwc91YFfQUXir3jTFSUvHPXwPu3KU/yJ1fm9rU2RDyxbxm68ao0ZZGc4SC3/Af6lqgNN3/
cYVGUmE8RBR8r4y4p9c0YBFcVEw58CjdPwzbTIoZM64avKl+rPENUr5t9OTDBZxMlqY1VuuBury4
/zLiSFd24qUZR4NdX6thPEXFF5Hd4VqdyWqp4i6EPYjMUb+eifDmxxE8pCBjLtTXrqViCY2OFwqv
VwigwmRaFfeVjOe74JAEMYeBaJ7AwadiJt6FWBuxp4eBxZXWmRdcRnfX3MaOokIHMe4q/8GUqTNy
8PIF938wd2g6C3e9nkbGyiEJyfT3fHqyKQVhtx8j7NoBeAXWQ6SuomO9p1OgRhW1mVLEooY21quk
xMikMb3JecvAmWAp5VznYcZL2hZvLIkydDn05VguSIZBpF4gE6PCALqxMy+LLxHsRU1Yo5SEaXsk
g3ei1ysX/rZGR+d5ty8OXfhVFx+BxAJi4I4h+jGhAOMskWlpoN0AcT3aInNu30UFfiMm+y1CACgo
tiWSNnShmfnQ1LlDhYRdGqLUSk/kA5olVFN9mJ7+LE7DOgtfjsc9OTfQdvS9VI72IOfqsS31SxLx
eu6rSATw8UlKTUb3K7xAT9p6xeLAIPdVSZaOvnAuofpdBrdWM7iqn8Hf3pdeW1y+IjR2CGp8CFdq
DZZc60GC2OKY/NMnwrFviqx/3jBb2GTWFGmRnP58l6ydoCMxqmzUsReA6jEabndQjTLhaB0GieM0
c89Lg1AKj3yPE5eQ+rH7MtLwp20nPvp+KlgtavpE7jFBgYdJwY8by+8PewPBvR0L3pguLp6/Y+5e
fqKOZjYRtvd3P4FAKFmNuz/o3ThjUcTce5AsdxBBiNy1hnNcntOdXT3izbXdzCwwv6NhnJqH6sig
LvLG9YGq+itEzERoRbcEMQnekUM0OIJzyZF6D6aJJVlvM6jozmr+F6KmTEVbdcpbljhaRLJ3ftvR
BzgWdo4sF/XnkiBpZBcPWlfX+WkZF2PbLQGNpcVPYT9HReC7aTkthrb1D1HQ7QHviv/od9scIzT+
Sv7FeLTUS7r/SRn8XwvT2tShJVv9KdcGGaKMcb0B/nIorrGN9ZlWw6Y1AEozbAKG+gn2bRNhJWAf
Uqo67hYxuQQboP0ZYizEXxJSN2TGWvFnYQNdaHJb/0oQROnVFCXC0Sn0YwdfVWAXKOWc8M+4xWHg
/9UbgBKZYsmrXu5aF8C9R7WMp4mzjyF1iKTJuT46GcrrYXsG5dTUYd/jMIq+pxcbB8d+Z4j/Mf76
D/+7eoJ74schIik1brwFsOjzWZu5i/jHLQNR9Q0ZpbsJhdJdaSO1gqhSblb+G0LlJhnyGc/IgoR0
jkQlyiHiZjcmq5SmXtjDNFYXcH5kTAqP6cnzikf+iz4HI8pok2wTIsnf6DUEHBUktGaUX9Is30Lv
bDrdGLT8Bgt9C8zFTws7sH7qFBTBgeC/OXM4AV1k8mqOdDs6A1k+EKb+kwXAhb1Et95dhZUjeXNj
n1Kqo5V1/JQ4VFnxA7OCPphL+lLTXgb+kv8X0mwR35dHu7XAgavPkRgetw7V74Q23t9+5Fqi12BC
P30rag5ENxNYbNVTH4fraWFidrneiRN0cmjSaiuIjp+OK+S/hsQr4W0QoFcd26tDjjiXNrNSV0sN
MTH9yjg8f8Y0QC2KYX5zFCpAp/gXHEzahipgOJEhys32uOrhMI3aUuKqBRu+tcFQA4dmmcikTlTx
8KxyZJTj3qwKzkHqa4ns2m3z+/0GMEdgGYfvl9QRwJ8cCAP2vAqU3ygWG3Y6uBKkOzbNhDD0KzqN
Ygs1YFsSvppIej1vbwlfozE6MwfMR15GMcFsFaE/VkVdn1HuMOQLFrTeWX5v6VGcqoXDqygWgdEW
HClYgCVCW+R96n8PwgSVzScG00WkBBaohjznIjD8qHWpB6gPuMOXsHrD68Pyo+znc0lLu3ON8r2V
QYZTj5u4X+z94eNMPbHS94b+8GDJ79CdL929wuoDlielrHsaDScahSKZ22ZC+8QvroIeeyf5Nq0G
6j+tlN/1Odjy6fWGs0JKOtOz+F5azouOuPqOOlOl4FHt3lq1EljAiLTAbqHS/1zam17/PyxZzJSJ
2E5LPwb0kogCMPgfERm5BmyRc3ybyg3HgVhTiZKwwaO0PyzlZYGZdZN567u9Q8Vuc24/+MhNoAWo
LYR86reI6wqCaTWqAYATIoE/UEfC/fqnDJLdXX2uE3HmHALIypP7Z19EaHh/0dzA+Nxj9MZj8qWv
OkOYQsF8jwm+OQb1xmgO3hIWU1KIOljoeu/jx2RuSradBq7bpvZFUBvZCq8lTYWMRvXZnB9b2KhP
pP/21S9xql0iqtNjnRkkRdMVQ6VSdPRsiM3FW1IpVNem3/uny3ABFYFL20TAIK/iNGBS0Xql98M2
qcgRpsimub4TGqOXYIFUfVZUNuYMz5skmL1YpRr2CWuk1Gs4SpAtFVzxWHEIN6xJ/XHC/62da/aT
zZEI3mbJhM9Su8wQahbeBUmucs+Tt+gViB8iT15FTiTqqGrxdHyYQVld6I/0SPKkNy4GBy7A1SMd
rLbc6bCKlb+tH1mVzjDHd/NlhPiCqPSMDofbsNZDzvgBpqZx2oxV0sFrRMCLZjaXZr3Wkuw6NUXA
nLo8WRm0eR0LJQy2dVf575mgZ4MPxqCcvzuMx4wMUpcMG1E5K5RLguB64Wm4NbNJ6H6moeXvi6OV
Yumt88a63apJHb3RlFIq5a+9QR5VXhtrM1IuAyRV385FA4uiCXWTn4iWwn4GryEYsioeNxvDKphK
3uKPt3Y+GPNi2MwGA2GIZ9ywf57xpAbEpVG2C9XnNhDOXFwuM6WdOZjyudgY5wYQm3tVk8E7aRBU
1n6cVQCS1zX3waCceVpUbtHfcgJx087uGNwHCg7wu1XbmXbJoZ0kPx8VbgWJg1fPlfvCrBVCTYlw
seVhNztOdE9NYSk/VQqMl/n0mOvd0kPZM1y/yk0rkaY4NoI679/VPTUdfLsThK4eBgcxPAfJDOUi
+IEqc5Qfv1ACwVfv63SKnlwujttD8Gl457X5yZyF5jKtr2iBb2QkhtCbVA0r5ofXXmJJlngqURuZ
3DuX8Xpsmoyn9DXoN9TuJIDg9FiG/RGCLImBWDndjWiIZ9bsl9HF3LrKkQd4RxuSL+4sKdUABorJ
9R3DLCyAcCRtQf3oM0WofzcAk875g/sgh8iulEpX6cN3olc9uyfecjwCh2uRnoIShSgizW86xfJF
WtVLRzbsqJu1CgnBe60bNdIhhfyPmzy9bhgTjn7VrV5SMQ1qrML79sQl6v8suqYy4lLflESj4ELT
n2/Sg6U7omqNgxVjRrbzqErlWlPCw4BqaPBNeLWsrqu3TEZ1gnrAYA/IxSTLF5dd4kB+8oSwlt/O
11vqwg+lh+6cbqTFfWolkkT2X4gdd99m0uGvHpKPcC0MH30VaKrSCLWlUIYeHU4Ah8diHCiPs69m
r9J5KkTqXuw2aqPQKTtlQlRgCJMUxsQUJ6bCZF4fMRAKScoBGaRvvvYaFPMa7nlhsCpGTu4hY35d
LDGPMCACSWM2Ov7M+Pxx9u0XcYczbmg79F8NXbS6BTi3nocu7jvTrPNLtZ9lxzhjfPQZlUUTWq0R
VNmscMV4uWp5UVMzTtpqT+F1UgTEDBl7x4+gJKLch7zeeFo6+6AOqRZJ6lmu1zDN/X2z/RMCqeSJ
jxr6hR9yoPVtLXU28MMnF/ASzy195qCjANVHznPCLjLp5UcsWBntuSIZdMi6LF3VZCT2qOZddR8s
OjOo7qyPujC8lAdl+za8kE1SlXXejNMYbJu1UOthXgbxtZN/W4D9+60t/xaRRd+544lJQyk9WWZm
Nax83tsdaLPtjNliLy79vvuzisr/GFtn2EDmbtZm10vquLW5GxPoGN++N9epCN6FJ2iwdCnlfQmE
1vQTbZ2k5CLdz4huZO6CGpZpH9bkIb93v44T7l3t9fvzlj06zNjqvln8xJehF2Sv0tNPvvNMe7Kv
uDgJf1B3lPoeOuu5uJybJV4jlrk+Xz/JUS6wradMHK9u4Er/EwWeEzcQmtwz3IUE2eKa9WeqlBNF
NPRnboB6EFvd0Yk2HyA9WBegJlhzmxiMfeMnwNaurVRsIYnBg/u4T8J3aVpvYZ4VnYAn7yQWGg6w
p1Z13txR8Cd6eFJsuOxaesIS0JKy6yndG4xBNL98awvnl4EGRTHk9yCWGMVdUt7OxU9Sr6cWEdnS
fL7KX/huEusHyeOWxjqbxJqFO7aJ6kc+PYnFM1gGP/FV9MEh0vpWqn5/Go72zFGrh08hyN/VUn66
TLqM6CyLjzBP6NIWIGtWwXvvZm9RIa97+bSuIB4AMmxf77PWPhApw5ZKCTGX4vV3cIwgSLXiTkdX
gE3Bdbgobf5+gjx/ub630gsglFUJtcE1I300jkPoGdk86K8cFIaxkEEEln9xPLb9eqGh0BuSxCY1
WX9LQ+HN6rn3a8Hk1fxgID4wvxzYjuh1pcTf1XBubARzLmhCBbB6yWdVDu8PcOGOPFaFnRcS/18c
Rvdcg/EARXGgPEz/M3obaD2CHfRCdVqb+ZSCLohGlYZ/VCbpm9Z2sjwSz04jZU9YAosiKQddMGvJ
SydKJNyxZ7xzr6L8FGzI4euhxgdrfmp72kThM+EFXT8A6iztTVNuECPwYpKiDT73jBwCb8AOLSwM
oLuJ3oQ8/s4e/JmDyzfWQuV15MiZsrQ6IYb3OfIBj2rYbJo24tmofCLRU7j6fD/pLWuGY/TZiV5K
TTiKOIhTqw6TkbBfEGUGLlkkbVgr8M2jevA9HLKHLrhU5OWD+sD11+3ReHVrQ1qGn5ekeU1hUqdC
nwuJMObvIT1GIVW3vqw/NBvR3kI6kqXTqNg+S3hS01LedvqFVWYBv1vP7DTFGL7sRX7J6A2YNFAS
ihT2jOeu1/UK034zMOkRnzOfuX0M5zuy99nLwsVMngDx/n7n7L57Ho+HopswfXVZeN7oK5oVvYJi
+TtdnpKw23jesUyB/Lat0oetVrlj4mRseuCiCwYYjXd4h+NTuAGo7giY3lyfdVhTqtZ+dnnpqfTn
eS4vxuF9IgQw/bZbXuu4K1lrhz2/wz/U5D76BqvPdDcDTIgMRuaVuuDJUMAm7aS65ruHimemSTI2
5wW++OrObZn92Ey+KcD++yJjeWrsZzLSUkgkywMvdUaTAF6BGBbneiLTFL8T1t0yIKhNStNy9elu
ST+z4JXtEndGSsVfobYWGQ7WTC/2U7u8g1InYI8UCXmBMyymMPYv/DfzGnxxtD7GRdxqbq2n9Gsk
DoxfMS8hqEFM/M60BMkQYUcnZtEKr3wqA7sARZfzbykLYCO588sIZCOxB6p8HB/EbnOxUdfMD734
TGYsrYAhlEizqaQl28eeKi6rjTcPDg2oEjGkWMpFG/wGRLP2BEn08akWLDY6NHIV2/BQYBQGcmTf
+oBn3h27iwHt2z2lFuksqMbWK2XLIkommzUfPx7qH4nbiInZQdAncAcK2WNnIGTZgwY/dbhKkB+z
eibc+IhkY2vUCaYlwzrgqCV9zXwV/qWYPxGh+ngRh32Fc/0SbMdYMR82nFgwpmtmpz0IFWbid//x
ZiYQi99Lg0rIKeyC1/+YCdZ8pSFsF5iRb85ivAbNYcO6vXIffHsm5Sozw2xk8zbp9+KQHCdOeEUp
qFbdUj3zRyaAyq6iZB4OcSTdfe97RV9TWWiaEn+XMugY6ea7/aZJLV/YgJlgFiuGl5ncLq+TGpWs
wH/ELLa8DWdAwN7cUZo+jl1Gv3lA7vriDml8ojcwAVcNiOd94OcmTxUDHdLs2bIEv8e2LL4f43NK
8TCIsCCXph0TgUCXaKY9MDnP0YUB0aN4u+Jw+4xFrSVbEQSLF+lS2ojAZNBokRMadxSAiRZ07cvz
oQ4mBQF6HYxhYBztsXnfpZoWxbTf7dT5LuID2xf756eCZlWxGOH7HLBJNJTci7oeKDcsOqi8eom6
M+POOXr0c3Gttazh+FmlhENEnCfS356PpYRG8KLyYWUM2XBKS4pLvuss8EmfuJmQNThxcryuhWTU
8xvttq6dAvGums9Rb9fM69jpY6HkjAo+2ge/5K9N/OKPt1uaVK1RvVIFUHoVrvehi2zdGBewVZ4T
F8iVR979loiZd0v9Idu3l3D72NAiVB/sj9py3E2h0i1lajfo8sXczjiKtvBmcpUCLIM7babHfZKN
3JBtsF3h66p/TlorwkeZ4Yq2Xb4mYJcr6cMKWgECz/6QPrvJk3ErntGOCL/3rt1/ZynToJhlKftI
1kY8lk5yh2mKDR8EYZiXgW59g+wEamY5A8WsTNl7EHvMWmj7RCi9REoR1Mz6TuSkfx+55Kr+Nvc8
Sn1WBFMV0bQwo9hmtY1H1SfF8wDqqD/Fp0wQN1IQ7Z5Pm0jKBfzjfFfERHkq1yPe6vw/Yy3z/zGE
2p4+lCTNbktZRTNcY0XD/xbP9oQXn6g9AIZDFI0Qlz7YgdGKJdUo1Hys28weZWM84ZCfOiknYJFv
A5eg46/FAkC80oWaMWArEvUbaNBX39VzYnp4+j7jMG7loFpPM3OeRJpulsMD379yDybvtR6q9F01
dCp1ChSWqYIjP5UVcslPCAfPj9tDbS+DRododJaoHlSz/RhSOu2/BUel/qknc6ZoTGu2vAYf+ExN
fm3oTr8M3/kpsyzx06Ir+g1ob2YipPmEa9iseNq8tDf2Kig+ngd56Bdxb7XKvH0PqZDZldASv/PU
bxxwBacabQB/SA1Lna67rF9WzQQrplRljtb4L1hjmayJeVmfFYG+C5JB6rA1NNAFw9JfrdFJAb3y
OiNudlJaAf4s/hMlOu+uOiLMNU9V/KkHk9rJmUvS+ccggN7Bia0SovRTI0DytaUFHoPBN3gzy1pC
34Ndbwt0Vzcf03Z1WSgArQu1KH4n6yos0vBHZoY8WZ6BlS7f7ywbcc65CHjKaNT6r2aktqCC6e5S
Ox9cSxKaF6aVEBs6S4+BEdFhvRvAhfEVWMlN7c8NF3vtLc1CN8jvLNHqJojWpIBqtymWJWk0r5mi
+jV3Yy7AhIZAi+DgcsdblAZMqBhFR+QaBKtCmuaVmK05CxJmnMiZFd972ivBl0uiPhGx52wE/ITL
ge3OMwh1tnmJnV1MNYw6zCfCx9qpQ0fW+OdqbcXSQbHM80kL54OM6Kb8sVR5FsBZSDsj2fXLKizU
B6fqEi+JQBBjOSY4aQpYSZbeWI9aop1KvK9Z48JXstJWsiWIzTtkJY3g3s27zWBX9Vj1T1IVyzUH
SFRJlGlR6ADq83c0fcljx7h2l4Ipf6vu8sVZiS+KI8ikrBqom9UvcbLacp+PrH4+vHe7646KFH/o
D9DkMjAr8t4kNOxZI/GDcBLpFqfeeDWanK1Y3SUQINM9HBg1hBRikys/oIjoC01dZcAVIAbomVMU
NVRd49YHUSIekuuzWPCmvRweYs4k1Rw/tVWziO7ndLhR2qqIat18G9KZCpfwpod/ufpOO7trNcxz
YJ5PPRm8heR0bqs9nEfBcO27A0x12NaDoxdTV820He7pIOL0qPJFStaggVOd+kzcyMh12c88FOUn
ndAHwWt3iR4thOwuRl2Mxqqc2SnQyUALNn0b+hnRaaM1Dt0IWkDjSD7RRyk5jpziwGvBl6Vcn9tE
jC7RlgaHmQENxCA+YfTnxpaVmKJW2zSZPx5yeDqUENdSmltcvKFSTKQjqOFCIWXbSFaZUQnU59aR
mhJwMDYV1V4K3QZGFPeOasZvYINDIhS8CQYg0R1nGk3fv5HrIS8isTFVgxYAHUmaLjF0s/f+dJGX
YPi4r0RwSwTdHBDqCwpe11BBC80KGLPmxAfZa9sr8HJSKOPrbCvFZ2Osnff154Le3EiyZ8o7JYvt
BosxTSlYTtgqwUgljAJpoRK997nNvufIFFjHaMMiRixl+Ot+9AO54fjNAT/HAcaHO9qpPVmbqI2p
y91D4+h8JNsJhJxYxB5tmMcvPuniBM39WSR2yuRAzjqPbBdyV5Ge1PIQLjSMdadiPUmdWn132dlF
Ptx6m275sfTeLoV+OUW9VNE76eTiby6mMxg/qc3H2vUgm0PWvEvvfTmWxsjZD9WAGuacak912ogl
Yh5+/0Vs/tMnsx1B9kes8tU4jnMeAinSfTlF4tZp6CFs1fEbBd6lhrQfRHgqCeX3RAYzn4I6RYNh
q4/EcGvKr0JPCxpWsHtyeoiF/laCHVKpVSxwfi5ZPb1FYGB95zr/3JOv2MAlYWeRmt3TBGxAVIrP
QfJpnM6R4G8rIjeM11Rs9cHlD7llnvatOkWiQ4WLLA2hDLNIJL9K66GDDVvguF1peCizA1TxWtpe
YiPkRSsI0tvvTQ+MOzn5VMIpYmuKToEkfDnxqgzQjdAfmf8+i70R9fWMkfC2JgNLHVv6izPl5fSH
KwpBoU86Q7Yu4gAUroNMNSWXX0okvOojZJ8jmWWinQG/fb1kSM9VuWtM7qLJ5ZrGxjKsT3sXn6dz
tjy27ZBNIxxcOHpMtnhiaDCMfkh7F5k6EDd7wtmoX4GJ4WWq8CnW3TEwcNnLFMMIisZ9AVV8+k9L
+McvFzCeiWAX5aUbmXHg8iSBPUXkiWaUFE9m842zjSs1z/XWJZRuW2+rM5HWge5GVfxgrMzKr7Yj
4xHr75nlcnpml2Rnk5h2PFpcSus3Axn8XEBSr0HfYsC4JNAR4otwGBM3DJy/6/V/gNggN6vUZZsL
Zj+DK+8jUDpYd+8w32JNWgnDUk8QrNU7FoR7h2Rllq/LuOl6SPW5f77IbkDyTmIr+DkMr2cONkA9
J6s4DcMGjWHfASre9pLN4TnUAigYKeZAEGc3hO+MZ2ID2yB8raj+eL7oPudWZu+zlCcfGMPY8XN0
mSpdBPBNdKhfqrKkPYCarwTFZ0J9ik9MPpVLeZtKY4zgGpD8jJOqrgbqYvM5A84A1r5iJS0Ys82I
D4nqE63j8toOF5SquhmlGp7dQyCOQbnE5VdoDuPifsQ98Uxt63uIi1Ik6+wZJ4iB7SXnGjBUR2QM
tpOQIvgE0iwd4GNEGE+HLyZQCF/u2iSRetY2KJlE7+YHZWfs90QPFRHSwM4MRPIUj1g2K2tKwRAR
o3/3dnWXQciKNtG0zIUoWoqE1EQJHEXHquHzeK2uyw0Vf+fhnoINjXId0KxtzcdZ5zzrpErAOfEm
d6VW2e6pogjSPQX9aJtmRU5ubgFLAlwh566q7PO8DaY32UrIoTXdV1dMdiSvaJj9n+nKTpk1d8ur
E1ldaVjTK+WDl/Cy5fvaOv8vrz8GvbdlAHe8487161BkTfNXbsc/uuMq/P+pS8gMPSczJ4v5YgqL
illvn1lPzWKDbnlTJJgRk0JJeCOE7xYlQDE0hFYyge7U9GDYQCwOzjWAjGi5K7aM/Z9mHR7aBjPg
ud2AzQTPx4HA7EOpMFUMgYKPr9ouMXvuAEoYwGTtIOdOcbLvy24ogWiKPwtlkpqlQTnz7bunhc6c
JIMLwL6KHrIXJnkznKr6W3gQdwOimaaqFxpByWUG08/hF16KMy8Na21B5BS++1hJUY+CEf7YLa7n
5HqFsb0hHAcUQ6gwro1Ma5unzygeJPRZ8Y+qm9U4sAEmzrlPpzA19oWsOlgO2xYXjWw2lGUiVlJb
gEKEnIa7I8zOzh7Vj7Jegq1Xd22EOJsX16vHW2ppqwFSWQIZWWC3iaMtLym1Q7A2WmL07Czey6vR
ZUlC2wdHShsNRQit0NmtnhcsSnTggB970/OyDA495ojsXpuKsqEFtJRtC7cDBO+V+5ruBPr5QSsy
lfe2bpQSauIxC4eCvXD4Xn1grIVjhjp8sc8itdp9z2RT9kK4Fr3igwsRWJ5K8j2hOYENTgIEbJ3t
s3Pq9f57+GQoJsUPyQ4GcmJ7/6WGZGdgi6dzqqbHP+8ugAbKsRV8o85KGRCaoE+sWHwqrrmQ9W8L
fDFFj+9f9ZV52vSL9tx56t6T0iT6ju/KO591n+5621A/QYzLe7dkeo1CRUslqoZdkA/DukMuamb/
riRL3vb+Mlx9QUNY+9+BlmAnCOEHKznPbGtKAXwukhiq4Peh580Q65adcB7KejINUaAdRgIZe3R2
WH/ZGn96/MG6GtNiLdnegqVFp1TGKd2GIZzIdMDp0CqKVkhe83Isy8xoR8TNM+IOrJeMgKVrBGgu
m/5zfj+oaoT+0P/Z/FapINdohIhWj92OO0dqNmg2oXQlLshYJl9+2ftvzBUpHeqXvMGZOnYpENhB
kaZRFZRPLW2xe/nNlWU4in9FgJGVqGzM4iUG8HybisTN6wCM04QP+3j2J0s+8+/JEZYc+S5ebxyg
+Hn4rXxbJ2WCO9Z75rRqbytbRNBmRxPG6VBr2Ibc2ROHwIDStx0klhRCj6+6xv8JFcfyVclliPWq
9sJsfiHBjHD7VDaPlsnKE8a04RQZGuoo7XkiEKmn1IpSoMoumUBc+VV3p0/ZzP1aIq3afh5VPgN4
23ISKwvlAdL7F67guUaEUE16Bn2d/cN9IAfKzKjFBpaH7fgENs/aAe3SHUZ22qrLYUi4+2BuZddS
jHLza3iZ5mWs6dVwI9mBy9FuOZe7iYFVMu6J2WyUZQ7Wy0U7hfc/UlGkPZqmwmTfdGYBl6wOSXJB
M6XE0L3vMb02Kf8wwI8LwbV1FuK28Dtr4ft4GP6LDCAfqwsNKBeSQcH/LfAe25HVtQHLyvyw01nL
IuaeI5AB0I+Ien6HZiMNUZ7Z6Tjd2yBvBNvU21bP3wqz1nd71JijWhzqYTe8spkoSg1lgshl4fG/
eelE6qckhVNfrhO8NOq3RzNAFaETjvhU0j9feBdRx9OrEul+rfLKNn/ZoHd8IUvp6v/3vMjT8KC1
dIQt6kQwXIaZ9Vmp/Jg621cwo8QbCSLyGbEVwnM+ffLeRkmZhbRy4n+b7tz6KOMjKdButRG8XPaF
h3DvtevdrV9wuQWrv963g8/YAqMyCE4ILNhOmpW1QaXKKm2NYb05wtLdxnPalI5aai6m5cOAwf3O
Fut2OZ4Tdrt370SffU0sIQ0bhw9Khn/4V6yglFrquS6mu+kxs4iU1AjbiRYgEP0gVIE74I8dk7oO
8gZsRew1JAN2T4Tk+uiacrRpfB5TGm70NGiEXQqzrrrWPlIam5FzJnIEF7WMWZAkVHAlsXshKIKq
rok74NHHjtfNvd/J1q5Ckz0WXFKN18mET75hAWjMMHC7L2lRXS6v81kWq3i6icFGjr0lXGgm72Qx
gL+CBW1rvVVG1NR3OA6piceE2NOvt1y1uZo//CZcSqvlWjk7ZyGftvA+1zFxenlVSlxC2Zisz/AF
aIgDItMEi1VG0C0EU9z88fR+7t6q+BoaVFB18lq7eDz+36NSCihiDQVVMP2QhXu8BxmynZ8YjUa4
EBSiqbRSqZFhjmdhwcQCFx2pr+mNOe9EQejeciJ8hbQ+HCrYsfdrkzapGJ5VHEeNnqkDZX5Lz2xw
Hz4yaxXoAnMcBOeMUdCFH31XA5jrmV3Xh6muCYFQU2KK3JlfW+XhmiKnxlf5EW9rVarRKpPPESR3
UehyvHnpkfkVPwTCTB6TIyngtQHB5HxlEvq/8pGrWmexTqST6gbtYTSKxYTNNitsOU+Tp3bvn6k3
cdY+fSBuJSYei8PJtvsWUphpzK6z/ZwOsMzrerGOfg/tbbyS+CYQD6q1aIORHipZ5dw5kZHFNQ0g
4W/cTYkY6v70nB24q6UqewsKPWAPfBeD0/vthSEARJV4hpo46Ztn5ernx2vMd8c+r7DcuhytUfaY
OeLee13j7THPsaG4Jk8i0nLVw2zxRidl5WBzd66ejNzAcxUJHjFaLAGDyFho1WraZ/y51LpvIEae
XkegvugR0xenxXhDxEESNC5nXc2fm5ISFYKINlffj88pGTIyXUW5Y5M6zrJLQPHK4mY7oMkMURZV
Y03FGddiEhssmyP+jEJQJvnMtXF95QHF6cMx6s/sOlcXJmKVJpq3peHWVJYGdlCMicqqFH1hnXY0
/yOXLaMZHLUO8br6T5yX6rNZOmk0VW90+qwMyN/WugugIxkFOg2qoX7GdytJ9Rsf9zoOg8tqft/N
myRgC1wsLwiq6pu+a9xwDkOeXju9pe93htizrHmXdC/E2kCRPwzwAgmFjZVA3gX7q41atgvSunfq
Gwd38b2ywKW5eexAjyWeS1e2rgctomkPHo1sdDD5Q7YfSFp/Cku+fQ1ffHW9lhSTf8CklJOH4ylu
dgl2UQJmEa0EN/vSBXDaCaj3pxnlIYZyFvjrUFalMNa8n0/hE1NOLuWdAFFYnescuOvKTWanJSNn
KJpEQ/Xex8w4glUAhu6KbTuSlSahoIzXWUJC1E9eYxHe4/3Y1vUvOyw7wjc+WTZJAqYJne4fAIT0
2cWO+uUzpWyPB2Bmchl0WmrbDNC1j4ydYBDUXfYeXgSxJLlSBJsBFmPtRxadV6ydPWh6k/VtgM8k
GcBXXBMYNaTqXgKjtqyQ5QgoBar7N5/KR0DcJxNpGe1Pxxcizs/c8VWr9rhvp1v7sGwvMa5UdY4S
f99QdG1FiuEMIzwJIMdD6RZ47Gevygq6LxmExwkgBbQzdlq090EmoMd2lfwwsTcVgbfWSDodGvRi
g06NzVreQGH74MhbSc2GmtYCYhc2AcW2z9Og3i8UZtHnMP3wrUxARt3HeV1Vu4Tg7iNt7qu8WXBg
059QZ89+KXmjEmwVAMWLwVlecXeWnUAF+b5wcFqW3E+f8bGNV19pC0/f2NhCY0nZXcfxEI4DOoUP
ED6pjBB3dyybMDyOJ5VrUP6z0qbe5kMYB3yHAMc6tpMvvlGzFyrmH+nVlwZqbwJFTJA5katJ4Daw
SSfGcYfr5W4sC+OuiRg3wfyT2DDRmR8shuJI584ra2LcH4Eb1+0De8b51y6TmluFdZtcx4Z7lb+n
ZtkiBlyoFpdO/o1MDwgz++e+fybIjEVmlmmjUWeqf2/o2PUqqcH4n95GR1a4qnzMaMRpRDHMw9Ds
71dFY6EZcdu+Kt3Vi2HmrHLFTuWHgntdbWfZAnpxKRQkndbIrLdPq1DlRLg6bCfQn6ZcULD652xw
L5U5B8ALJlaOVsoAkEvIZi/opHyxTyYp8yxXq30JqDIpb4cDJMYwLJP9nHjuKwYyVd80Wnv4q01M
/E/QM7IkU4t2/RYRjGgULAPwtl9pxm/m5X89o1Y5T6KjZEgGO6ct8nHbmfEDox4sylbOY5FWn1FM
kb5Bipt8KsD63kh+wWrz1RH9giz9qvcwKedkzKAShaTHhcT5AZ03Qkgl5tfG0tnvZS5xPSJcuTXN
67wAgMCMLaaV8dKwM7OjFEEWWy1IBf93WdCdnxZlA+jnSRpzWCHvpMlEeg4jjl+LTzz0cMAaXBPG
6/SlV5N3KnLO1mC71OXo41uYVY3YDjR0881B4aDYAP1Lx4y40zUjW8P3pRk3nMjcf+9SIrlaIGxF
Zm8Js1V7XwV1V9C4TpyfjTbKVGKicaeyqH7tZKM3nNDere2wgcquq+f8y146O6NFWLYBJ31rW+/D
Kx0uldmNnD7eaHsIHiOHWtpf4QRz7oAQ74hLGGDDCiJih6891axRg/S6r2i77Eul1H1Kr1oSYlDR
IgZNn7pv+D1YhEXdVaTr++YSPGIsS8BRqjAfeKECmlispvh19ekFu/qRtUJWnjc6VTSrL4higf9S
1c9A8ereHdGjxkADyZVor9GAqzf/aK/r2V5387jUi9r3f7WJhnE9KyyRuor4aqC/efjmYDBhZo1U
mitQOaaee4NvTJ9+0w1MRnTqWe5fGrkXsxMv85JDjMFdZHWb6oT8CD6MJHRM9sMBWgMuDCUy4VTD
4L/e/VUZw8znIINb89nSMTwNucy9i+cuDDzvLhFvMbdTlzoLW1q3vLdUfPbcxgRTma6x2S41jjb+
wjqWfdi4NiqDMP3xhU1STzy/Q09GxPZ3LXOZbqKCrZqbvKXMmQjsKz8xLtLGsNV89XDIryvo/Oqf
c3Igliu+53c0NmnYefuf4aVHRmkuOG3sfugl7Ld38vkWlZyBRc0rB2Lew87lmd/XZGOBDQHBmfzk
1vxMNJnnFNXdRT2BrPwetiWtqPUTbqd4eS9XYYfPMJJSfKdhutkXAqk6jmie/A99T3k3sTsHOH3B
r3YrjYNFH+lxqFsKnt2+Y2csH4k8DJ9l6HsjZsWyQkspnjdo3tCdPpcJiXYRDdSHrOB9nAd1l85L
ZiHWM+A2NoPzJYn7TyKQZClEFjsdAK6H0UpwQpqxjhrmX5WTzXSoTsY5szfPyRS52d/quQGccGZB
Qk/Bq0afEKz/R8gTaVsIWGZPpN0Wzscv/0IoVp/EP7pl6teZVzONRDkPu6Z/lhOnt5npDlmfpgUO
u2B4SUp3ZvlH+2GcOHRDUQ/0S4zNhAQFwj6tngSFS2eTHVnDCJmVDBrbhXIiOIx4nJzVVjSD8pd1
1TaVsPjyvsCXQFt94uH3MTpCISGWjRiC8AVP8zzRiirfjeG8CU7nDj0Tu3NmSRlIOImfbV1ksSah
MBdMqvwBm24tkK0ea0q/EmBkvyqmzzVaFU25fiDAtP/LzkiCmE7M+xUpCwcZPtZsvXe9yIxpYFkQ
Vi2vV7cbJjjigui7GzLI+NE0TNQ4r+/cGbeZYQqoi3HiKsm9ef/P0Ab7wh+p32mc9aFwQ6S8NRJ9
H13pKN+eXuzxb4mJY6ZFHWPw+ssGAgCslfU8p4Lxlw84P7Guua2F4repPsbyeAShSq7D8lJppbkp
bWXXUDl0dsBiLGY2bKkrq7nUsI+GjnxyCAt3IH6O0NHG4I8FKv3IaXXme0+iWnR/5yTai2T2x8v3
y5ZRBW3HpbLWSzsSA9zSSFcHKwZqEXCXo81yFYQOSTq2sglsWGUyfCu3s/LaqjIKE48QnNAad+RB
rDAINictLM8or+QphDDP2Rm8mOf5hm5IV7p4av3EGzMfu0S4yk0cmujZMYveHmKbo0l34kp7a5zO
36v7w+HHsZB85euqcoVDz0bmxsisMgnbdPJvyrF8BLHsWZd27mDuO2xukc9BEuoz8VG2hqGtKE/9
eBipkZjpN34edQDLotmwGtB/nq3fPAS0vet96rQlkELRpzHl97TDvImH3yVs6/sESLk6X8LxVvdJ
a2KHp1aYYQlDEm7+OnZza7C/wV5bh+AWUd7DygYKksiI50jMEfbJAb0AZm8Sh80tIDygRwrvIGPY
ijsIyHElWApVJ1onHa7qnD5YnEstdDGEbq0K2bUWZin9pln441gDk/zIql+xWRajfYlzJtJrvoVl
CgENKWU3zzGoUVxozt/p0XPqUlNf+YlTpS/l2oenLMa7vgKFOhMoLsi/Me4wcQPtDpjF3ytbD4A/
xU/aF0ySj5xz43YQq7Kr1kpEX3V8XOX5IkLIoqEI8sFYWtSK0mcPuUK7/MWAmPDEZF5xELKHvTKe
RzNZe1K+mJH7Aw+i7Ojcr22TpvzAsWsWSDFMtuxleHE0h7Dkwvw7GE6k2/AlmjDzNHVQ41XNSvtn
AI37xK3Wl00NBY3JrElZfMhJfERX/y4bThG7w+/QjTKmw27A2HIIjTRBh69LAn352soRg7n8YqVq
2TF8v75wGyRjcH7hx5A+QdZKqNPzsZmjc5DLCYxzDo8lAfSS815vKTZZes3Zi5n5D5htnufMh095
tUuFcoZ1OIJN+iEayMt7eoTKYg6mFfr5x4VZd2BMNixtTYmJzqt2IACm7th+++NJVYKKkzu8z8ET
HvGPmW40ceyZyhrNgo7Lpl81q1tLJqUrgyKZ8ruyDCahj8iYbbSoeYWy7zpbZpajShGyaGwC2nWc
l9mHY8ZJOGMVOkncgnXWm5keMWIxOzXuYfmlDvSTp7djtcm9f7eSzkmEgoHYCwtGOpVqvShTz8tB
S/9QmMZn4RGaAl2qQCdXrsszD5BkjhBDiqrCsp3LFk+tqDgGIPunP+gZeHmDCIDSKCTb6ukhV/10
3Kh/V84v0uguDC0ulyQx0fYZ76ypIEXh4T0r6XPxG/pKtOkm1wPi3Ur9jsfoGdvwfYCDRR4n51Tq
LfKX826kPhkN9GiLr+rsiMxmatYtuU1Hi6PKby5X1JkWw9FsW6L19FJmqQhVyFMx03n7bqY5+CqI
0DLvqwg/9/L7eeHh6t9cSEyK1QCGjstetBMxPIBf/uTiipXG+YzMKY/D2flAewCCH5USUrHvfmMe
692KILPpgo1QwVZo5pHKPsItxENDqvpVReMFJjGBQIW3fC+Uba8nRhHqiag5Oxpgh4yZSGqeEz3Q
Q5lCaNqSYWv46/L1YsHWRtfdS9n1UBGE1Q9NY8TzfhYej1JMsuJyH9+riO6XEMp66hxTzC1LbM/E
kgH4SuPqFVco74rHU5mb9t2fH0KOASxJ5r1Lyd2SAPUTwdYoBA67TIo0pdgrg03ZzOBBfdAOkY8B
mbYwOs9oX1ACezD9l8ZUTg2Ux7QO0A1m5E0onuWc/chWaEU4GiVlDTRqFdR/s7qX24pWurGYyuyV
SdMHQSHicYywjkQsPf9uy49rwAS3KZDxHHk68tKJ/XxwhniSomm35ufsXCKfU2FpafeZw7jYw0Ki
wW/Ai+mUrfcCARsLBywgzxdWmv2hvQsbnVPq1OpDVjcJjTVVTTtcDfXGZ5weolEiisubnLNTRDL+
uyp9c89pZSlQd7SXHggBZi3XS+Z5WilkrAOgof/a422NcK8oo16H+niKSOtXgzVdYCYshl2FgToS
WsBDOgWag+ZpMbDBww5gW6iNU4dYoaV6yKTEkgc8idbMhfcY4BlA+fEHQ8kRCQKShbEt5VMIjOGg
a6RWZCJDk4xP/MVICXr5tCCzkIl+8l1tHBMjs9bZBpFftj43OMwJngoJQlDU47XA6uztv1tTNazE
64Vt2H68tpaBOicN4T0KEpZEOR6iNdcHeWTo0Pxmcl4Ka6JohorJCajSEsxEKDyLBJjMmt1IZFl1
zgtBdaEpLvZbksvhENqXqaQYpOoI/b7Kh3+vq6BPSF0kct5/NxSKwLAZ3ibGEdNBgd35B7eu5Bye
MiyRPsVzcCFWggYMM2mMjitFVICN1yOw/HiM9PHKtQ37akKAzno+hTJH/EpyTa1lveJaUvh2GjRt
clA+eQV5DygRUvnHW8GbHrulSYH+U8UIr79zxnHb+jWySmvwqr1SCsxqSlMttRSiA7JwfvIIWeB4
n8k8roOTXo6Zq+aPmdBDAQkKZtmFJ0twpd71ShbjiSiBysvTKiPA2EqypaCE128m02W0gwt82qxh
XVAHV04OWgoBhfYSs+5hDRN98kDcfezBec4uoYNeouX0a8icj+obFBdD07OhQVBr7tmYFXKmQplc
QAV+N27cmHyOCBzy1Dfr1iLqUIZGqam7G+p0KN/ImrTL/nEn9Pa6fmcIBbmxVl9+GAEddlJgOi7G
YNPy0PGGrV5GLRs/WEb62kixGmqN0Ec4ZhCgRwcMuYEkVbXyxb02O9eW4rN9qzInGRPzE+3q0vro
1jj+sgeJKQwuIHTm9+rMVfOLkkR+tCl/TZA6AtuTNkSeim8lVZqBgb4kMnU6ZHpYmKb94YDV6d8f
rrXO0kRxhJ3+IzNYSJxF3zpsYfZPMlikI+q3MtoznfMg16/9TXUnH7ad7W8JmdJKAx6gCWP9ttYr
STa9YzQ6uS3/ZDmD1ms9VMfj0hBGv+v9CMZjro4EN7K3zGSzwgxwAR0GXQj577Bt794bu4Qy5Bqc
hraJzmC6yMuwaTTTO+r9wSGN0gTF/aQoVPpxcJHcWRKmb9fdvVXc8LB+ra7p4MI/UneABGUQZ1Hu
Qf3aDpWokfzRLZ55YHeyJ3CuytA4vuIUZOdLq1cYl/uXuAB6HR3VQHUAZDqYyDAi9u+4NtRDsLaO
6FxlEBvLHVdYc7ZiEPSCfwVm77s2ePcv+x9fw2k3BI2mn0+ncWJc396pIdbBKl5f0FoHkTBRZxi6
ew8pldpWGbdTCYj5J3J+7DTMR2jnTlSCDah9qXmhy2Lcs17EBZkRHh8YwqFXHzBrsSPpgxmGzMlz
DIu4SKC1Ik2OU5hHjEDlB7BVDLry2UyfuYAt4DWiK2U1//DPvMc+XGWkNWQZLEYKaAuwa3GreIEC
ouHmQCwbD0Ra6GvFRFwu31G0afY/3pj6BK7zti2HRTm6GfN9v7NwojId0fD6WZbW5RuWOgQ0z7nc
uB4Db83ko4oQmFoV2cQBM3/+XJrTEAjXP8OBkj99hWBDG0CkF3TeUwzU5T4gjlc967PQD0vxI4/H
pfbj/lEGWRppNp4HB8bHdwAOC9MO5t71MKQD7UXwlrvnhxdBlbbzbEAtg6e6DJuK3QsFxoYDH8Bn
fGHioYXkpSvIfka1F4xBMjFUj3w9e2g/arR6jDsEEGWHf4IyoPygPx9K+rHMy2U+WZGZ4gEAJ4Sl
ZA19TbtJrUwb4v49r0TbS5XFIZeoLAV8+PSBorWiC2ClEmb0C2QzCNdn8kqPEpouoIq3kADpsUhp
iIUccaIoQMPaUi7oVjzaC63FUK1+OrKOx85CXYcdUb5ZPX71nk16gMb9SYbA1xFRIizLR7DvC92j
lDWIjp3MnHdeCNeHHzvSaZsWC37Da1ht+ggnaIFW7qeqvagyCkPSCoD8SyaLrbChCWDP3GsXzJox
nN2zT6+tHd0O/K1PkyNxkkZRfCAWLoxXSNrDBeEN3R79Eb/rQJXmaQqOdMOE0VMhyq/b25smB+/F
f3V7xiV5audtuzzXLkI6AuISgLuYpre6FYKpAUH2C5kE9gDbUwz4HCyvT7bqCr6vQH22aq3A9NHD
+OBvF0spT/CrkrZ3I/gK6mFxSf6ZQKFRVFllg/MkM1mF+fZ9bjpUoSI/iPv20ccTOaPzOyG1upMT
d+zle3ghZbzrdDGIKje4/+oK8mkkQSRV1oEg66LqexgcEN3sPkHYng5uNUpYYJtScGUvBG+6uSPn
dFcU2VfYNZcHXvh+2w2N46BTDHWlmp22ojmSrvMMPRTl7wxii12Q8Wddjou0ww7ew7IcdmE8aQfd
0N6wr4vFfgmZMKGkNotDAiC0HcKvY1jV5J6jLmnb1JjGA6TNjUPGvXWp8eqZNBFUoHv9mHt8eMPD
rQ9b+aQlRIrefDFADOs2LFCMlYAiFXAB5CPUii9PO5Kcbsl32V8XHq0WQofkXN2ZSxiew0CJKxo4
/5qMkJVMsfI4GmSvkNpRKRdR6vpJAUcL1SrVlmnFqjvRtWpE8a/1e5UVhKNUai6mjgM4o2V4FN59
UbmMtq06sNobel5V5EKGIUsPiAFX3+V9v83/LttrUKxV/T1aZsJyDEwriPFZPkCVmr4A2rdHrzqo
LKGt3jt6G0VaO6/GwH8Xx5rvu1cFPsuKfew/LjDuVtAMVDaK4RWvH8mUx4AuSLZ2CbeCzBVT5l35
1AhmMQHBVP+gjY/7rzL9mtFHtq+8nc1JXzTc+goencYUrxDxsfCnvgu82yUKir1Ot62fqFMNDIoz
Z6f6CaOSJOitT+ajfXLt8YFAQDnsbWjm86OvxFH3q4SgCZGaMVhpc2iVbOnTwG/CeglgRCup3iPa
D+uklQqMU4NXYFOjoJFyq5b7K6tqfbPKInBKer7DdIaxZz+h7BjL9PsVTJ7TeO4g4KEFyNU/U23o
8+3h7RiJlp5pvrNGf3i8q4ci6NY0VoQXwhw1dal8D+FrezxH6oa8K3uhK9eMYJ6l3JvpMll3xmb/
wsR/RboNfKfW4mDVGInBnDTfRTR6TzvgmTUQ7ggFINGKWtd/O1nC+wEFsj5ztY+M937KGZy0jrNq
snrJ/FgDozZ+0tX/XFwUEt4fEQ5PphBNM8HALKbiRKoAfKORDkrfQcv4IkqY6sXxfsMjCap9GLPd
u+FDzXoDLw3sMKpGdCPzc6MQpKpVnfVxjvLWvzsX76MevRJ54dU52u+aKD//3OhdSCIroIpMU7V9
D60GhhU5ZfsnD2AnZdP0ZlcHGwhPD0l93TWwlQD0a2LivkL6uUfwU1RQiOvqwbg2Qs3h8XgwoUsX
bR0wgKEI3isrtoKj5kPzgF2EmAToL6308PyEbnIiLNZXDdf2ybJl706Ze1W0F6PGelgc8L6x7T1x
cg1kCEurWzlU/53fvRpcGxk5C5fn4s8SfFNb4imOmjb/V2naHh7U3boYdfC6aeFRmnVrOLOz2YE2
hq4vxmrq8ZjAIP7HqdSERBPHZc7GQhE38KstgPI/ZCoYaQCU0hQabiazkTHvHFj6ZxG6Xo8zcqO0
lH5VeZvb6NMS1pjpQySBPq/JkIiSjTkFsYy3jawao+YVEhJRBcYIABNKrj1Z5Btxu9eEmrr6dxAw
guSiCYOp5hmZNGDDyndYm1a/pnBPUqdsmjyY4ohGVgOt18kTrEUdpOsl9B7uKqY1Csjy1lEzXVW7
ZwT6G2IebCX/jr6O9XXlFL1dNtTw2gSLdMFa2pCHm82FZLhdbKeK0yhygyKc5aYxvaX1/KdAalE5
dyp3pIhzTEiV71ao9w8LQNIdYKSENBBNcVvNGL3XDPrkQhwi4A667YtWVEQOfNoIgUqWlcgQzA9L
rpGcCN2nI/GT92srT44pgS6/lxhTp9KiTC8D3rJvnp4blCW2RnQrzXYfHndqv6TGGg+2qg4vQRFR
EhdZ680Pp1BJlVl876VLVWU5RNxLHvvrZt1oggCpr0PLoiKc1gV2tQ+F9tM0pyRSEaXug6BRp6jW
eIPuo5XvS90lZPkpmWSCw2zwmb2M0pFqyBFm2jcv/+R4oJ2jO3Ft0Oqoy9kTqZ1in73julhRIWMh
qXHtAlrJCur3xLE7IaPxYVqb1+9TPLoRhwniNXKindDTXqc8mxzpZZLBb+pGMOB1eaXW2OwB4Lpq
kT+qzxMPBMy41foOb69ct+/CKaKihm1SWbyIgkb1kGQ73kp44cfATucPBqt5UBHU2Ntrf7PEiTQr
5IEaRCQhx4hGSk1fdHcgxHbdRi2VFcyyBo0HOeSBGcmdppayY1/DhlfOMH/Ez/UvFd9E+zZHCieS
3wbUHxGpWXd9kq1yQ9r13oyFEM0ykBRuh4/NsrgSWE2bsmPzyH+dzLuagS/dEm+C+h188bpSVOs4
WYZR/cJJ4FX4NTW/s4qk4DdJHhrQckw0OfJ9DBn/EZDhnnT4gb2+0fCkQ1XV5sOGNH47iN5KdDFT
Hr+paV1K9xpYAwEWD8BBDiZ43PClgUtUI9l9VE70LWGv5tzmJcK/WTGdQBQy0soJbKNHGXBkj45z
QL5y77zoWusfPB9XQnV1Y64txlcm7u5DkjWyxtbWv0KgS9C4FZFSi4HxAN64kLT1ZjYMCm+D4s4w
NX/TUmjinWbJREYSqemqKY14H+x/TEiD6jVjg2b++TQ8woGw1RarYm1YvJyEA3XTbV44zDlIB19C
V20prqF27vOYMht0ncFavsFmrPLSKg4jHJ8UjBxcKoReT2NZH3SBvBrZ2P3SV0Iuh07ua8zpc3al
XX4l/hox7N18ky0aBPzl5d7XbF3OA9xhl58vyw8U2EvaYZo6Z567d4GEcvTt/PhbP4x8RGJBk01y
Y9DV5fC1ghlEzQxI0YF5TIElms47/+u99UO9hK8jKNj+qN8dujCF8ztWWB/uqQHKd5b8I656bY/4
fXTfA/eeWNJo7xovBNIY5tcmggHSHXJ7S2+z3HdunvEKp0+A5+VyomszvEkPecBHLE8jAy1JjgrU
4yIPi64GRXD22rpnLi8q2lmzq5Aj+BMmuYcBocWzOJF0mrGe1MEk6cn/I/qmEhiyMdJ2cnBnMHzh
umV6Zx5dkVQAQvGAyJUon2W496DQ5BTHWP0dVPUi7VonDSvZ1J9EgRC5VROh1cgBsvh4vOYtt7yl
u0pRKiNRvSEGszNhjfPjmlUnIhQ3se030nRJgs9DWGtZcdUNYtmJAXs8KC31tok71ET54JjCyKNq
bkzFzZefpFoBnXeCJTGghkgSt+uOktBlq3C+nm4GmgH2azdvL2d52H+FUllEhRe8qICpBGLBlo+3
hCqHYYPitKNUfqQL5Ku1DFuuSzqbGT+tKdz8MtlWgCmVANBDfcJkBFd11Zx/mZlJLbGu346+Vou+
/urneOZDgTDtARNPPYshkgBo9wI+gGngkdX3WVWjNXAHSYGHfTky4/LQF/qn4u6Ydl7M3ldLwY8M
sgdv1s+7OW0RNQgj0sUi6+u8/4mU2BUWHlzpJzKL3lGqGmS02IbmbOfCDtrTQ8fuWywkmt2i/ppS
yQBdDiu5QK99xi8kBTPBfmt3K4Ier5U29Z5+nv4DrZYpwkJH4D0EMKeIS5z9+LvY5btDGLUuE4+7
oVnP8tZYQaNSaeAWWwEfcHw2jsO+t3aQSICPPtpVDJ1jj5d9Ue4nMYsOMDp+CoLWLBqw3lbRLMse
Ok1ug+YR0Eou1gWrAUkYFW4Kar3bvr3E3Pttk8vXc9E8Q+9bxQshF3b5qZ+n49gMwX3kHpkEM6c8
Oc86U0E6ZjcxrjDUFkGJSvkkpp5bHpzemUFD0KEawVactUvVXsavkliKICZbJUIFFQi6iVVhAMd/
3wqeKJOgBgumDI/K5xz/UAVa0hiL551gxYc52chbWkQAr4IQEEtfr9NPrYP8MajRJRtWFiGVIdbZ
/uOnTiYd3EvvnjpDcMOAzugTgtGL8uI4cz1RU5cfmz4+pW95d775bXU/TAv2PPaV5W6IKlMmGJbV
Wod+cf7ulJrIh0KI89xssAcaR/5t+Sgl58vhDYW9wGmWjhnq2Bd54Mw8KuULRB0GP4jRnObm66K8
bO4DXsEDLUkQ9uoByxganAcvxRO0w3e8I164R7b8KkhxYjTAaMRhS4A9Ojy4V2LI3Tr14WnG56iS
p+mqO4GP014QcmR19j/qbiQD+VMjRWkFdli1FspwikrhD1J50lwBlY3h+ImdlY3DC6o8xub3S7z9
44khx1M+dXO+aK9QnmF0pH3LxgmTkhUIJGY7YX5rX2Sx9IH2MxGC4CKIPiBfDipCteVOuUfVKir4
2vTDzfk07JNkt5UblrlDMS+IPsb/q23ZmNJSSj1DwexC0HCEBxWrjKMyGkA0UuikDVNiCO//9pw+
EaZpobtHS7mhhDbUfEm6IvPobxMqi/QzGx3c83c8ayq785RjcAmo/TbcXJMZo19awE7NH2+N7wFw
/SHGrc0G/dEq4Bq6UWO/jBfzw02xJtB+XdiDroXtFxvohojuR8lz95Dihfb8PVL+B9UGlKpHxCO5
0hHpjLgvJX8HFVHdp2ZcJ/gmfZu4qU29XYzRsVm5S+M0xdZfQB/3145iYpDTRnCi8jDD6hZVYbdA
juQWfK07hJzZEvGjxsuNG6tlsCOBdYScJg5BhRb6NB5FSyKLw+NUwpNxJYT0SNcVxaq3w/Z8A/kW
ss91cXGKlcFfzt+33Tv8IlDPxaQ+UjlOrJCq5UoIUD09FgPV9maIr0BJ6rjB82PknF+4dpDYE7v4
lhjhrqVOvtHMhtibajUH4ZG0be7gFjiNRlemDYUv9OG6RBEtJKvDPCL5PEgm7gxKpZC6BliPFBMc
VeoeUXH1d4kKwXDqDRFAcS8JClWzz53bcaNhB8nbXRVyoJTuxM544r32M8udHkiuNiqgP1nY8m05
gR1iKzMV4iyYIQ5qu3XMwQfj5t6WPpgEOKkz/+g/sr2FEH92plax7Sy2G5umbiyplvmX6Bs/8p0Q
YpqvA7Or7x63iJ2Z9DT8TdRFjR8oX1iuiTtxY/bxr3vjicSra/DNTBA+8MdXDaTgk6PMbjvesXyH
imxykTHiop+E+PzqvatPsJMkSIP6VNueYXYpOwWUf5D7AL+uhdFGrjXoBdJt7ND/mtUmDmHLRGHg
OPqV6Pw8hP5jNrBzgYU+Qn+8XKix0YyawJTsbadtzTwrul5n3F6t+DTf8EUZ14uBxaDrTf+si6Zl
BMriPXYLXwtDyAXjCtMVeUScwTRAWtiQ8YHx0pCTjrizaj3Lz1GHwOKmeGOclOmLsqdjMycx9YNY
wo/GoSVW3DHVw3KqzqBa/iSwDCJKIPmJhJdXq40Q9/yy/RjMY0ceg9HSQiOrjk+wOzbDbPleVWlh
t9MVXsOfpa4SA7t5LsnYvOjld0noz7MiYMbNcMkRFKFAM5AU3vhIjKr1tmJmmlQHDSwyN/Q5A+Tp
OFbj1wvXL/VX5LyHalXu3Mi+zDePGp0cbowjc/u/5xujBol9X/0E1RQmESN5eua27DIjC/tdvYOB
kh9i6n9tWX6+DdYwGoHdGjCRnFRbSO44uofx/jhnE9J6w2zrtInqCEHAoi7XrJ37NQwj3+UFASnN
bBf2SB2rv2TgPDBGobyYNPGbPpIcybdtKW50XCtnDdTCv3LAzbEkF7NcA/oK7VQ4blYqu741XqMs
BjJlZmNW9Y25lbwHrRdxjCylCtUKw3ABZaUih0j5Ug+chSyiG869nq7ye8z3np0DP39rVsGP4PXf
cUtrmrh9FE6RtNq64FriWu8nj/1EgE6PPFx0hselVRH3pilWILu4YTSh5mX3U2PxlvPp8LpcG6sc
7GwKca55rOlVKm/CXSexRABHdzKfMCbUqdLNAaIAsKHTSjt7Sy0luPw30OfqVjuxNtWuuAAgY9ll
FnUsDPXuTNKAbJ8MNOlXKHKSm550ikyASrujcO1Wy/IPRxBvq9L64PD4HZ+Cs6iy4FVrf+Wad4VJ
opaAPnPYE72BZUzpDJzVSP89a7st9A9EKKs3YfA7KgFLoeZ7FUt3OpeZjFMpR6AgdNa7RgsFxodm
f/+vxkSAQb+WoBXczw4sJnCGgZl28PJyFEKQPZdeJfQvm30t6UuNvpIamACIs1YkMP8ahUfTSx7g
vUqfeRZXbIxkTGoPJCdEsR7PVr3yL1UYT6haxDf5Y19jp9NG2D2ZEbWBvX5FZ5vvaG3sXKK9q7yZ
CKAiIoa8T3TkKJATD74TU61V0j9HMnt5gIPllgHS/ZuJMWVZgDouBuM1yK0mNHCGDrbiOBP0csUr
SBLIC1M1VZ9GbLV1xFs/Kor05Xl37SH8bC7Uid4I7V3lBuTG8iitj+lbmnuZPyMcp3d+ut38J318
BvW0GYwrVjRU+ChgOeVlGVPEsuVSdbVnZQ+v/kK1KtvV5LQ2D/pxg5KKxQ/1M0BOgQZIdeLbvWzk
3FApaGU42HDKjFcIVJ347nXjnJlG53Zz67tJ2wz2tmNx+kJoB8vpRmRcRygkZe9PNgvZWoDhhVdC
zPeFvIumHMdx6X0V0imV76+Zxb9+j2HymK4RhMngx7LZOG76WXILz73kXi8N7V+kJoZSulhgFxpF
RzlnktxQ1G0qaRbrLGHg/XIAnfq1DNiJfmo1NAfbX2hI201xkzR6gWpBv8VGp6q7mKBbAvmIsUaH
ZjSutkffIiPnAd+s14tbCT3LQWJQF5ZtaHLG0HFMENcZNEp1uYqIC9PUWU3iYfOwwd3E4IhkCjRv
WqZMDdnKlYQ3o6DqqIAjamTHvABEPODVW4ufkrRQyXuOURT4YgEYf2d/iPSe7m1EhsPx6bE5gyue
3xhUsizj4whf942NkqBwvmTsTqKuZ+Z9Or83/zX7QS4yiCNbzQA0x60/x+t4Bt8CHvrHHiOnr7aH
zBkcjeMbotqHi/VaqIjv98lsSDD2zmoYwRsGUlGDZmTnMlz7KEhnZQULLJuCcdVXBblhy2WKOs+y
EMtn8ddTfcKkhiSDcKp7j8Lll8w4G9/+H2tOb+XWkdonUPRJBEAI2KHCJNq6VKEW7x8WF0/cEPEj
bVXvce9ji5rZNs0NeOarRsKvB3YZMChK06Qg8ySTJttwUaUlRSsHT7plRq33Yvwn6/jZRFfcwJsR
QI6HWAoMEFsHUCg7Ze2UUo6AcIo9ZSE4gmAXHtH5v1eQl5fCPFLamoAsZ1D0gax3qqfXsxTYiVoq
FbFSfA1DGkb0xdH/bsBoFabTR8MBrt5kXFgL47uQEC7G9XjsFq8pXaY8uGYqYzBhxv7Kqw8X7r2n
t2zmHYOfbF8+alQqwdZQF04HG2hTqXOXKOEmZiQlvpnzph6NeYF22k4lcOYVPTWZYNcUMmT52iOE
ExOSadukl9xtpvgJpknSbcWErEhSgA/qmCw1geDYC7b9A2b065kpqIwJLW2upXzpygN9vGxo8TcS
Zd6drD+4JDBnaUVL/T6nd7j9efpvttvTVwR0iaHtakAHYKm+/40fxh6OE3OXXg4oAQqzTDJntfNX
3rofsBw0/xoHnQAgUcnJgVDXl+QHmYLT+4iOFhAlVvAsuzxxzUOEMvec5i0NIoUH3e00Mk7YqelV
zubc6jHkahewO8Xbjrz7/b87/kIfnez09SH9vK3xsuLQQCPt+iDTvBoRrWC70CACIr7UPHoMPtud
4s9c3+GcMVYrqwRAPG+30PHLmAfoLpTXeJa8tdv8Yl5KOaNHzPFDJPlAHqGumgQ6UHmO+HmewF0u
90XvU272xt86z9ZbntgX1dw621l18TXnihcVFKnoOXgPGmkp7MJCvHa4Fbvbg0GoiR3cUmdgBJRb
0ZlbHaqYR7TshPWegp/1WqNJ74OH7ioTXtyKXXD78uJ8JPkQtBigmMex1NAnaMsLNaJ5L2mZyCKg
R8fiJyAuv0BnvQ8ZT+e7wlN54iERhjbq+lv9ucGEL52FHrNP8FIYXYtE0UfNPel4zeNLAPSccOjN
cojDPmO3ebMiVpERIKMSL9rQ/JeuGqzeEOWIUhxdN8s43JSDHkHoQ4T2Co/EHzxW8+TX20ewUQxk
PZwF6LxvS7FIOR0RCqWg96sUdIGUTKgiLIyH5MN+4CWUIDbDLI+Rt64eKsUQz1xZKwaxZwDyqb2x
B5zD7zqNHOeFYtdd4gl0Uqh2cegORO+43l9NYkZ/omK0Y3LPbInRDc/vKvF6/xvUHCB4gw3wb51D
/IvogW3PWGF2Xc/WZczR6iWtM1fvRwRmgIejTEK5Lmf/kVXUENIp4+S3eRAsUiHkcMH6Lna8/90j
ACQ4d3ZuIPDVUSg7KeTRVld5937Z/sJouSGdvZDJIIyEjq42ABmu3LF7za/PInpb2wXdoqcuvyuo
gYUhOPIc78ufBFopStQHCFHL2zU5W4EryN2vXkvLLVsV3hh82CRgxaop6Ba3TzU7d9X49UOBNnBF
A8PkEIqIzMbkw7dLgs7lEqkVSBzApcJb2A0um72KeL1ejnv58zvhVo1phuAzKjP4FqdwWLE4nKhq
UpXa8RoxkxNMPUninxobYYbOJXFhA0utYiJe099ESoAkh5CrinGzbkgJqjUGjX6vwpI3R4JPFA7H
w1q83Q9Lh5aTC2YKD0NusaLVuoEoZqUFejomqRjuaplzXDj39bFKNv8115C7bYofYF+Xdy56eJso
a0XRJO+unF9Dc8Wp+t56Ma45MUb2tjBmeS2MohnsNUfN/9Xu+yVRtp3xH/8ACtTlzoHBLFWYfrUh
LS4iAmVvVm3OZT6NdXyN5pBcTkq54zKSqiD0log3uIWr6xu2Ixzf4mdfss8qz/ZB1AbHhDUOE/RV
1yWplKNp/CLUuXK2viFk/MYq9YDey3TX0O8iXhZeAVj9BxW5qW7mZRSsy0CNmd9PrPPtIMGRIBtw
NOK9HnWNv+WaIRQFDLfX7N0sjHgG4YtYXuCEs2JycvFpsjxbmoMlHvbQhlZ531dVcjV2ZMxSaXQ0
SbDN0/NhaEfdXmLcrIY0+IktNvfoipmjtIgk81mPGdA2RCVqxT/MqSBz3vQPLcYkrFan1JS7+PGQ
CtbdsAF0WvVoNcQtoazxoO2nRMk3WupFEi5D57KngT0ruqVS7ZwMg9qoE/cei3TLVqa/p0cQLbt8
FfnMg8EpZSVx1X18iBYoY3X2gNILGeXNvL2QG5XErzhudD06XH7P3DtJKI7NreBbxDehzf6Qo73s
EL5uZQBuzhT9+ApakBvAJkv5jqCxnD+FFzRMYsB88W424b80aha/V0G2g6XmmbKFteS5fb+9qRGa
uhHVpSRBOfEApZfyPmnUkOGUWynGdhOwRuXSCQpOCZmEhnLCE1i3J8uacQMwg++Mack+4PHXhUlo
olvg70nx/3hGjWKcEYGHmHd9tBi1hWBW57dvQPaG2nm9YJXBeXwUIUdi8hYh2xUAm8O1QS/pR6xZ
RsOtqnZcQ87p5/Jjkv2FX6j4mRKpyrAt9rF2WyeukJXZcW/ERKo9NVL/FgikM31I4jP2YV2ThOQW
kv4+KLCqa/YCtFneTdB/QdWbmUhPcPNALxU90P82MYe4bT/9H0WzyoPrbPo1M7TeLiNH8AKWBsh0
PvA3XXXpNBw78ek+bIVNzPLralbTBVD1v/Ob7dKc8q8i9jm4WgaQaAqGndnuvXCM1G1/x/ikFR/0
ITLpj7k9wH7a8n51OeY0I45scWI5TcIXfm2iEpuWrmp015MB5TZRBxDpj99gkdh2ANAQHp7PF71V
/eXsQ3l8qRCgZrwMB1EV+em3CONmHfU6xItspvGNrPWSDMv5ZHc1luZ2HmXmGnhQskPETvs7+i3h
yb7pp5ZeU/FBnEkEVKYqoN6Ls8AwAvx3Fn9DRY5JiC/0XRMASFZl4lZN4fZ9Zh5bz6Cfbyfp/TsZ
o0SAOz2gCSUFc+OwHS/5sP0pnu6RbqbP/IDN14xubMzjHq3IEuwnFaHSGquUkHrIg/kxKhWnVdn3
+piIKAmwLwfmLpDAcw3NQOqQWQKFz5pimfJDX4JuuEDSNO2NnUCgTDrkY/UW2vuNhN64y4KGNERd
5UpIF1cqvGGL6mvxUK4ZyJ71sRTqy2oVfmIjISmIkTGxy8UlQAmATZTrYtrqPckHq00ibFNSW9Py
0GwOVEIOsCzJU8BWxYHLkNeXhf23hOcH7cUQ1VZfMHom/TQ8LMWe4zQlOHej2IR/+WpPGnjkpcTD
82gwisTiUhaxenN8R2lseBe+bCb4GeT6e1XZsNC+PLxWdCeJxRk3tfJZJE3O9rtnCSSdA/KpVO6B
nz19y2f0wQUI4nLFi/Gh8W1gSUULgN3snaC6xMWCSQgAe5GMN31yLdp7yL6pdVntaJHBESB1Vhfu
W2PtzG3IcQNm0KKr5Qvfm1lB2vfl2Z0VBA2f9DHRbWyNLKftN3PAMyll4AjMWsjzlefYG5xNIMC3
Ltx14TxYExTs2LlZtdz5oKZGr/BlzJHHfO2WB7o5UI0j7OZHxu3CL0+SSqycyEBy7g56IeyumkUd
KF7xOD/K4Me7Zg2EZYxSy+Prdq9+3dOiB7xC8gHsVixBaFdQt5xK2ERJaTU8UMelgB0ni60Wwm4J
/kX09Te/zPuOMoTkOPsP8MBbQNkxIrpkGzPwj5HinPuNMqvEoAutgw1qsNDuVexyFgHnasg2cY2J
U59/zsdMdyJ0haj19Q+L/AvnFlBRFoe2++d+Ztl4DoJoJSziUJK0q6Osvu42W8i3CCcnpk/kzP4R
1dYfII7lsyE99rOCgl6SRJFiXeN5uXSDY5Wd4GrccVFUpmsIHiF3YI7c0gFrO9J0XcKin16HqUFF
6gBqiDLQMMLKUIqf81nvnLnj7wWl/mIRp2TAhH29Pe547kZMj0zavT/S25xho3qd7r8oFL5Qn1cN
F3tHL56P7x/nLtoKA81vi2OXRQxHUZDZmgnHj4jnahphA6fpq6e4ypl4OFEaTJjR4vYXk6YXU4YU
6lj4P6SqD9gCDJTim1j0a3tB+pJpdmlEgwdAJLIEl70fEq/rnNSH24nZfnTrkiEyu2WHNrNdfilF
rUdWqsA7GKc3NTLgoxrazwa8PuJLpXctWfbGzSlDmfkUV9jdRgtm2d0D5sotzGYVsXk+ooHK088m
IFlYBcX17ZtxhXDbtGbZqrZBZFFwu1NnhG2Ekb/VuyOeu3wzet5gysEoeyRHvBFg+PfsbKeTm/A4
32iX/pDrHu690WsqdXZM3rTH3Ozo4pPc+b0vwyRO7odE31mbztiv6IhvH4Ws/+TbO1ZX2hl8VfFT
LM/LZeD7FqyyD3huicJso584n63JoNPvdDO97AQOr54S8yPvQMjTwajIvAW9kOo6KCKfb48ntKnf
ia4vyw5Kq8kXuMuK55zig4qKx3uuUQkeLoy37FjFcEEQcDTuKUjrq+wEnQy04aG6ty+1tsvW4STM
2HhrO9pMJpUnlZukjR7BWlYy0TWGPOcO0An7UM5xE9G65Kp1/DHSXdDo/drrsrjchQlqXM5i4P/w
fr5oG7uWgXKuaeT4zCO+9I6I2EGJrdMp9TcEhmX2JKS5bxHT8sJqZkIJDAu+3s9RjSLOoYFM2dhJ
dddBk6lKm2rAdLMhwaunYGbybEWITUXaOyQrO6ZluOQHaLariDAaQ3nFJ5WqgX/z09ImN9D91Yo3
h8WUsNbYFazcE/4q79bO/aPu+1dJSBQomuGxbA4hnEaTMYUxK8lhEvawDFFb8z6tyTswYFjAbzV6
/zl9AEc7G2vyoaxZuUCIX5YeohfAHhss2QD528taql1wCiXVjpLulpJpMs/vWFr/bvjSE0vfKLxd
bt9w900UXXlEjRfxiZ/MNqTpiKdXiSIXuceL/CyHXT7+RlcBnmC2tFapL7c8E57rChaZxZ3N7MP2
Q8mjNzm8u1RbMmhATU9PbXMIJsza3YHRlSjCheMqH4XE8gGPK2gikEDeYhTTNFOhD7BwhQzNgC+G
aYkVeUBZitHSAthUsWR9yGkW+LlYLd1YjqBBReUDEZsd3/cPpR4WejJglnVXZnLC3slN+8CliKKh
d4tT3dE7AEgzhgq2MLntPbCDW/5v4WTR1+GpQj4RluETg/5breEX9PSD0qnvVwiAgEdJXCHKGAPE
b16rgROrfKbvvytfL8LOEf7ChiiuDCbskA1w4vxm/5UHb1MC7bUfUptXf6pLedSQE/ys0iML+2Wa
kIkozLfTk7mG46Avzg9QJwTaMvGi6EAFJH9jID0ne+glLPTahVbOC2PU8cYdWqSBy0ccRMjgNp1o
n+t3j9lRviFoN51F4PYJbcaEWr/WPjdu3jnxy56YXBoABHCWUHuJQZ47Ixb/4EhqBBdVDFa6M0Ye
h+rfUtDODF2xtlr+3VtgxAmx6rmtY2ZGuzR+bttvs7Eud7W7I+/iCjvgiDS3wEgcpZK56DtLee2k
WEY9c6b11u1jBQfcGPSqctks6sD0sHTpI/9JaL5LwxlRWHFjwZSYBF/QzEZIK6t1GUzN9hV8Zc3m
byNBXxjwUrAuRdyQ0dUP4nJ3wJGxkrAhja3hm9hn4boVY9b1Jsc7q7/xyh2XUk1cpE6o+V1//FrV
ba7TQR6RTsFU4rg5e0k78/dPLk0OvEunp+6nFacMiAWOmwV5k/ySDUpn+egPtcFWYilxfnXY9p9a
AsGzXcUYHqStx+mm8JqUJ1ncU+QNh3to4tW+uj+uAaThcS69Vk2yzXD303FVbV2D6mglq+R6/d0A
Ytj9AolTMZ4XAZ1FtbOwCtHW2DM6adV6LrSHhgOU50l7F4kn2zSRmo7mNNCPqx00WtLt/6Sj3Iyf
+wSJeYWtVTsohpu5ctoTer4LC+BdrNG2oYDtDZ17BDv8dZk+KVxp/2iAzNG94ukFLfibE13pfyvY
F/9WBBrmcDH6eYQrOq8d7hnXLPWaLr0DUWOVDWt2wzJuQsl02jQqgPu0XEA7TCS4uhMsSs3kWCrq
vMowrGjbo0Y3eeVIs3VcWL0MMlOp4BK2+z/8kBET8XNKKLnEudVdF3ZG4vI3OZKvLFsiUArTJmTC
L+Q+r55jsbtB2lrnPIVb8tVMsIyLpS7X7G4tpYhXxbvo/53frTB5nYWzorhD8HnLl1876JlwV7Pn
/zHtuhvMFwQ4wLive8s0os3n4GZaev51lRGVKZNBtV2KWmelLz/LhuWv9AI9MOb80yKQYEHh+hkA
BNCxLYYd9hiUekzgOKWj9moJzZ7DMo57a+gC5lAGePbFAezDXG7hyUAemlzIUf5UADomN9KXGB+1
KlMepPJmSYb3K+zH4pXwzl8OxFmHxn/WNCXteUzyl1PDiPwx4ddYVMNNeiuog4BlSUZiFQLBgIAQ
Hvvcah3lBjdpM6g/DEc2T/vXQiA93bccr+/945ng/td52Rpldq9ZIBRRneZN4kVU3xTpbxNQGfzJ
5kTczUUMGujAneB/fsx//Yyq4FeJHBjSHQxeO7nIrkTBAOuJjtNEn6nBok9UMnRd2C3Pu/Q1j32l
nBbG7aYyi0GW9YH7yI+l3ONI29Cyd/ie7/QzuG/I/JlwKKsCjQVtD8mf9bFnm9g/nNw2v+lrwO7x
m/5wHt2HcEN+QGmqKNBUT0YpsdR1WdlR4UFRD7qzNTI2xlApy24+xub6z9XANl5kdzFn22b7qFz4
MVmWaH9whB7SXZM130OBBeM3LhlkSeIrHOPDULN/flBVe5kT9my6DE6/oD0yKoAY836pHvmO3aU5
tgoVasmtFnOQME7pMCnILCTi6NIAoXTtoJwDf43s/HBgnZWCovZcCdzqFvrNgnXxzWm3uPZWRM5y
spbPqG81QyiHq3/IxiauZy7TcMiopTA/oylhc0OaT69TspPLZ0ucEWJlmn0qcclAqCDN6l9QzoZN
A03yaDuBm4aKYxR4B7zV/ZmdY45VD5lQIWhWkfSSghedU1X6Q7FYXcdrtBf2ziPkYwxOWhi/n78y
TCaLSAMLp3UPlHzpPgyY0/Qkk6DJyWt1HjJn7so4/o3mxcv26gI8dH0e22xwSba1b+0BCHn8AJls
3tgykvcEj9rUosuaaQv67wBdYYCA3nGlXtDQ1W7bJfRWo3ftoaic55kfQBL7gudom/8rpJ26kMam
rvnJ1tNjY5OqLo2jVN+CwVBTZ4Z1OTcsrpZBMvkdfOJ/CXSG0PW5Omg11W5kgd3xsOjnkWETtGft
QHKoZeFqA0U5V31lweaEavv1WWciXI9w69Fo2PCk51S2+a4fH0zMvkvpXoLmLFAA+DAlxQQ1YpIm
bog5fREap9EC58RQDsxCMtCSqsOgqDQpSAolSi5XGiMvWln3OPqgGglQol8crWuNBIpxBX4MMxhX
Kd7fBBycR1+HWEHN1qUoAGSEih0mL1ZBASRg4c2pdma06OB8sGXrxDhpBx6ZBecB11TJnelIM/iS
Q089fxhDAYMTfVpAcE0sNckpB6tWLz5Uae3vhCghHnJVE+oaVvcKYD7XrX6xCSwHD3hjtCM1opDF
lDelTGrmzp8+xr1hHy0PXVJ9x2RaQk2JENer9G4cjLUO/qWf124pIBs9IjdTOpeuuFZVIeEKWE3M
qFtfFa348Pif76FnzT8DAB/UX7RYSGWyaAsxw+dyl+JnZz7bHadSvOK4Tb3LvSR4iVnBlf/21/K+
tmbAKUo6+InbSb8uGaiqFtwUWehmgkJ9Je5L6q2TwPv4gZN7xrP1im75VEWO90VNnHccOvaO5uDb
3ht/pDU0WMfuMxjhUiwuSac3Ep5ya97e5xJG68JUeTHe9OUpHM3BPqoyN4n5I2u6CdNUa4h+EMrK
WqEvxS6Xc+pX0sqkOjgBlF8tKdDTM1qpn2jqIkwbjOLjnZI9F2FuMLe9ElUyITBit3Eo9SPLyKvj
7O4322QO/06vbWNt/UOx0a1iDFhlm6vVi7glt6cYm+vCQvZw297iv6xc1W9xrfb61cLQLCkmqJQX
0SUXxr4SC1rJG5Yk+61TXZ72bMoO9E7m3S2fJXMlaO8YTXHS5vzTupnExgKvW8EVovlfed5/tM9e
BKqoWkFuNidBIxJ4/LZzDs5bASAtMx6eck+uEsXSaNl2uAFjYzQyWaLv+/8TvloMT6PjdmdfE6B+
NXpQ69XK35dgQ+USeAitT7qgYIZIomzty6Px50mDv0U4CmxPZSRpkFniBs2LwQwoR7drAYWD1342
Cb2FxbVR85uDLYeoqyqHIl1GIkI0DoPHmThmL9t40Nw6CcJXKP1h+3C+ALVIRG1wAZcvlh4NBp++
Ii9juMoXCveLuSjx/4LiQP8jGrYJI2JtYcVIWau3oVUfl66gt2+LZYY2yfqm7pkXqp0W53tFV33h
f8WwmN+5vBSOIWjgLS7VEhhlFEs7aYrnFCToyQGBohHwSOMn4eeRvREvOy4Mo0GWc2w1IiKh1oCW
npRb0AbO3FdmElbSTs/Cy1ZOJYuieW7znBbxrL2s71tTCCkrmZt4Xklc2tuBvLcO84HtSA48jmEx
wyTE8nxEPlMaKf+e1p/W3eS+YK0NzIwwJ6MtHcLI7cett4BfbrwKw0110P8U/ll8CmIryU48tjGN
GfTzAI4Ey5clNpgmKqJn6zRg+wgXf38Wk77ThViESRltnEKHspeXG6I0SgrFMef2wlQZWlUVcZez
qQzVlcQEvDjOaXYe9DPi81m9e4u3UZ8VN4kjoDYlNhEU7of2Du0oEtRInaa9kEZ4ziR3M+5R0VBo
mhYj0MYl7pgdGOvIDk7IUdOsey1mUlBu0764f0VfPJ/43dPfUQp09eleoWlynY+IAamJanFtQb64
ojf9TVPaFT4x7sQs55bxFtxTQzz5tAhER8BVy2p7FxSQ/0TAfznR9QKdcajT5zM5HjOIDqME8Hk2
X8oPDsv3sUsy4QWFaQQ+9cpyvKDdfySAfNF2EQNS6KxlE9mrmqtf4630OU8UXZykN1IspYQqAi89
LeKzIqPxO/TCLtqLimR+OFvdY1VTLskY0paNJ5n0dPh+QZLgAzln+q0SJ1X+Zex7izEQSlkhrMD1
Smn+kZyc546Ll5rJRw1lXlqoo29xgBZMmGAgEQWHWFSIIB3drYOpMsQB0pm5MdEAjG7Z9Mv26w0z
igAM4ksJOji5PImXL9FHYJDF8rKC4eapCb8b2uN5EZcO9kEYIf8kDp53mrDkbXwtA0uMtZEZoGs9
18xfFK/PeEqlsR9EZAdkLdWg8/5lGsfQ814jMB1/Fe+AO8rTVoyDGvB0XdSrAw6EpuKNw5MiGhB1
3aSFPQfrJ8RYXXpPmyq3P4bzM1m1M/cwPOcIhZddkrB3SBTZEfcmcvomQUvN6C66ZH3mB8OmLh9A
0VcfwPTRLf6GvuLCjl0vpe3A9YMTtxTouWZB6LM+M948XAiEpJNcIvcVajn1uX1dBm+lGsXE8xkH
hhuGXc8raIi0dl3NWjbFJNrPGXRi5F7p9m84IDrRBsrnWAK2VPh7LSbuATLyKms26Jul++wR9Bm1
KiUttDHJJJK1EBv2xaSA35xaUZ4ldxRR3ikdpQo2TYiZhOxBX1ecuwTsPMQS5XgLEiveUydQ/nL8
g9lU8WYYrlPwr0/TjD/UjcH6u9Q/x0WGd47f4I5K7JvycgSUzQYwo1dK8qhiyX83ubWKTMKMvwje
TNMFdrPjIq+O5k+wWNCpfXhVm3YMZihc8g/VJKBf4OSr3Ntxlog8jOTQOi2TlHM+MzTZIa4VHaob
XYgmQgAI6xlpEpwp7+J6A9vujU1rQtiyB3cbCDHM/znzr3m5p4D6kCQgHZpEERzU0tqOn2VMRLAw
kRe9Qxq8o7u9ob/EofMU1qyT3xl0g7EsORymxpjT3CYDXGIgIug1CL30UarYiG0501SZEpIluZFf
tFZ8fDaiQ5BJY59lt85XCVZWT/PDoj+Jnd8GFOUCNk7mWMRgxIKmkX/JMXN9Yp+BuX1WsPE+As28
LRhKgVrHHSb+toaTQG78NBhteID5HY8BVdc+SdbVF7fRGC6c4JdL42MDt53dC9BkbyN9ilGxGP7E
8KrRPDahnKXvhtTrYObZd1DL1/ZP22QmsZjA0/LBqhOC/NY58BFXaSkB0yBg+U2kW6A/YdOz2vvz
JKJ0rO47IWM1eZ/FCGfCiyNz98nItZI0QMbfcZhclUOLYFf4nyPXUBzohgAHzQR3f+wJXa28thw4
4B8kdZ9g4J2Iui1i65LNxMIxTj0jtz3+fCvPOcte8qdZWQ774eFqCz/Ea4a6A6lcdv2wpzUu8rTs
bB6IiK+S6f35iy0q2JEB2IEDLGcr92Tx9vV0AMlFT7aaPukVatmac+ZxsASibUDbJ3DI4RpOlBzS
56APl/g3i2ufFZWxgC6MLVtCtkThuf6L4JLVaiNMc5YEH3v20y7q4h0er3b7fE+8IJntz6ynms0y
+5ZS1Xo1VxsHJPJBPRbEQ9KvtvYMCVmZPjZjeQLUUJ/jbnQHpbtedNNy7Zp8uVMv75iCF4UjoTBN
moc+ZK7nMv/tTJ5Z1oWA/2kBkeQmHWmQ8p7VgRoHOjcyAlsg4JKkb0lCLyblNFypDEpMGhD6y9ip
5UPyMmHhbs6FcBw+5l8QiD2e5ghTrXsCTqzPvrjcZOKoX79lmpFzQbUp42VXD5BfPtQ02HxeqKA7
502/ow5iVGkge0JubDCNux/aahFIOv9NONwg3819lmrWoVeXUpeJF5A73gAFBHA7v/sk7PZ8IRcb
oom6SxQJ4RDGwrFlhe+beuSfPSIh30fsUo5aLknEevGDA17VVIclPSV1WspJa4/ixXG4775JpxdG
NlfagZKgeEYECf41TXNIvK+TcFaN6bsfPH26AjcoSEGCwgh//kKkujMjMqCepYzOZ7uxxp11W+O5
e+tPyJymtJfQPcmFivgzSxiCYJdAqGSoeVbKzYdeRKkCnzKbGb7nEa1OOa0x/Ocy34GQj9qgohrO
t0TvpedhPEY8lxwORV4SXXM/fAh16xsqc5Qbbv2AhFOwkXjAglQQbgOQaEfmxtfB5IjuswyBE6r9
RPlzYsKvGvolV8OLipMhcDIrvankwtQ5EL3+H0C+RYpqfB+QdWJCcUSJvfhah4KsoPzZCHC1b72n
MblRl3qPr9UxzM2m10KPg/L7okd9/v2Ic11nnRqKoI+hRo2kB0lv622TUvwLf22bqU8nOoSZAPki
QrEX5iBiLgJGGkQUnEkUOLrp/d7taMk0xp6J7siOtErMIT2GIkhYKNIVlxd+PT2rro0mg5aacH08
vDMEgdaAQI/z9mCZ5PstAhI77igL8V4GJrwPizkGKl6m/yQl/qwK7uGPLAoWUaJb9hGMgELunhW6
1Bzkn6FmBjfSgYcK+k97AUeeeODtTPoC12zp9JAdRMvsOIXEat4dOYwVu1f8/Kxyangbs3YZYKhq
yJSIMflBtWS4+ds4URDnZ7G1kGyKpcBUL/xzXFwAR43WUYa9apmJMn6NqNh6a/GtboPK5fUxmoou
zWzahlZn0JcuZYVyx6T0DGAaL1rUBnDL3t/OEdu34axS/hFeFFd8kZUx56TNricmBUAJK502rjL+
eAM1ULIvuf93HqXvCAtji75IYPw8AooBeoe4HdaypR4ucPy6QLnIzSG8DS4KS4PQz7K9h957GfiC
QyXcD5mBP7i6W91TLKs64zhNxjZ8UO3g/r+Yo3dv8QOas5MJFjGBfOP/5kUCouInarr5HqnEUuX8
aso6i/CVUPMuxV7zOUTljzMd1IlY3mE1LjjDxF2OQFSBy75BckKYmM3rXJr2m7hCfeMQXrkOsPzB
r2kbwN3p/No/IM+dQP+b+51pz2mkDH9jWMAUuB50TzuNrJzZxXYXHYBn9ZiLvaHkJJBuFM6At9YB
tNerAYcqxOszCJaBzQQ+DlcOpRy5P8NqqcE98UTwYeqUXSt6l5jZ1rkfdUKr09zDZNJOE/ghUC9m
VvqJH9/iN3xYRQhOiqP3HEC6jEyqsaV4G4zUCqczKzYJxF85gd/w3zTr4lRFZNx+hudz4b5ImSCl
Sd5qJQg4L7HIb64WjtXnk3Ex/dA4DgwzQxK9KcRNULI4/ZRAixkOzGJlzVF3LklGgxdpTznt74eI
KzTymELCSVJzQB5GIhQ3xV6Luq112tbXNnS+SH8xQOe7x02de81ZHOD/SahMyLHiTuJXy402VoAx
ZYteiVPygQIIzw/LY4EbHeQT7y+fDPOBRf/6YscudQjovFvTUE4F5niB7m8MA57qWQ+A77iMIBes
eK6Qwh8DGavKX8I+nTjqOPgZC5k2ZbBa8tkBFOHL26VN7wh5kbQoOTuCul0JcdM06M7ZK/EmbEKK
x/FHZkUPrdsJAV34RZqLyxFCEIRiNeOrkDM1yNmkPSPnKvvFlw1kaVJuVPAk7iOt0OfTS8RScg38
EcKDVYRu+wQFulwEO3aRXHYU9gG26NlY40wwqu0lkTnNFnV9DMEtI2wP8/SiN/koQcSKcVogX3Uf
ouHsToSyodr1qSOC8LClZY/qKwevjII/n8Z3lwzZBs4JnSYL/MD4dlYmRVuq/C3RbuJj/JK0FDKx
psVATc4p7IA5oPqLoSeUV2apGiLMjCfAEkTgkOj3PAi4aztrd7aitcDIDRsRkXsxgQD8N8PMAbAx
a5CPPoUDM6/POX9MwC+E8uAzIDKOtxgukNxTSqab0hbixHxxg3/Rogtwyt7HzeGGkl8kXMOrSQL2
CYLRpuq26MF3uLMtedqKWzLVTlkAOhxDI3KVKNMK+mmZ88vImlCW178iev+0CqXi4n5bbgfUgg/1
ILt55Dbf9HS2soV7knNb8CouzS+UP1E+LNrkl/9ME6Rx8Cc9I/DKxzoEyW5ohWviwvLXjNUZxCbc
I8FcJaszEnGzmErCIVlWN33Mz7PjO7BJt+IUsaGzM6lL6WvoGQ7HezlR5XpeCYP0iLFYSWS3mjKN
JUlfM+lGS60YU5O9VCbqhbPS9C0A+eVCeblUeHVbTVfRlCDjyxqnCzrMpYdm3pcd2JnQBL9d39Dy
RuhFr1xdVd1G6bOcQszYmhV0rGghcsI7CvQqupK752vIwAfLrRFHwBaSsNucz8DqaLSq+tgYsu17
LSd3aMdFXaVlDI7QTB/ddE8mTRbSGkoBuTDTRoA3Aus8zwlONYp56AI/5zK2vOH16Qs4pCTf3mdg
ZWia4e10TEFN3MgsBKTAFsX43zyKU7Tq3eGafT1UzdnPrhq4SLzc6FtpXC0nqJUwkAmRC0mfjBU7
Vq+zGTcOXCZb0nNO0Rauwzh8mOjX+VHU+dmMg9OOSslOi8D0kTeG3XllNYaWk7CqkarzOz03E1UF
S16bch93iIj6LMdyeMtolm8H74joGbj6TJi6fO3Gvvch/hMtr0WSqYtx7RMjb883NtJNrbsWCYl9
ZYLEuq+80MyWo7FnIGBYMVsSvN1aSkaQM2Z2gjVz7XoLmUXN5x1OmGov17PoeUiWrI2dSl6PZJ9+
xUhUDlLi2nAHr1hfYWHJ4UTmtUq0B+S2g8r24E5ui9Gu7JjZlCZE4qLoJhmunTn4Gxzg7LLRHdOY
cdSEcKe2Y8Dqh4PUWtzAoGgOTW5zgBqg/J2ARkBfVy8pVpNHNkuYJDX4xRC9haP+2uamMrZGwt/x
sE65Ts0vEczkicDveXABy5e8zq+G3Iz2tDUqNQW+rop/QeaA7BFbKM/HVi2gu73wL4eeBVgfzfQa
GGVhBxtkMpujKyi+u/iqLJGSrZEympXkSs9ysYo9/BHH7GDcSuKj13kb9YLrj9fmW1PUUD/lrWQd
DPUCevGTssMZLHeoB8X+22EtyqilMtgJ7Cxnq8Sxw6shASOn6AOj0jPwKOzb6EQGxlfU8LqDfac/
f+YvMZgX2Bo5tYAP/UPyuCpFsPPsspk2WdXuMz/4ohO7jGUa/eYOpSS1TNA03JxLCdlLnC3nMROJ
QFjj2PDHKP+/LDRxrGyME0jHb/MM+byHL6oEJ2EyYNA5bJAtlPfEDBqFxB1jpXpp8D5MAYdmWhiZ
V/s+D5kIHDa24ge8nBt3IjzWorXICYUT0L84elJB/qlRaKuW3KEuSmAp4+MIqKoOJIKkHnCEzSbm
4oAjPKpgK90c7xTUy3/ykUNVqXu79c/8KH4CkyEAp41rPTz+I3rPRxoo6idDSCQa+pssL/uA4Y7Z
X4XT+gu1Bl+BygRokMIug/qZ3zfYNz9ONbC0YJBpr0IbIT07r8281yFIjj+Skjf0B413isk9BFpv
q5eE74SO59fwuYsm6y5JltOj5kosG+2bn9jHasiyE3xXN44J3gnsp/G7RDXOiXLIF34Br/4SFC9z
i5YfF7V/XJan1RhfAuDLEWGRa9IiJC7XZKm9884rWXTFnY60AeOW6GEfyHwWEbfSqcjjXHqLOahX
9MFpSDa8ff3kjjsLOUMBjoDfCY10PtzqtSMzPYCL5h9lMuhBWGGXXqTp6cqVJpQtzHwzR36OPt6d
iJEeyjHYiNMSiHUA+OiIdH2JAAXEWCfOYSjONk6ZQ6EzYBUlDxpyqfKUJogLjWLaFYcYsDLGWvTg
tOQHfN/t5wcZXGfZMF8YLytcH58nERouP9N6xxuo3V5ZNHGVdo+4CyF9hn+6bN/ixBiQ/KFteXW8
gKn9zOPjNXC6oXWf6hSdYWXzttSv6u0fVbY5CLa+3Q+WjYHGxZgF7uzSxsOzdQIwRhtizU6FdA7+
R5CCFguLacBrs8A1OPgEprokYwDdsN9FcEO4tyhABe3pFBSzVwHPHc0YBsUji7BAcW790zZSHuir
ZOODvfrx3PBp0oMf/ApPJftfBdyp5q2PlQcWset56Eztl2iokWcHVRfIuFwEPdhub5UxtYxvL2My
c3t5ThrK0Xr0TygaCKdMe8jdYwgd9MDU9Lilwk67LIK4JRmjSA/L8BsIhOKxXcOS5PvoJrSNgnnH
secidEmDBjn9Naf9WcpS4JV2z/AIy9MjyOsnAWHmPpLkwwrRE4xBVCIx2UdJg6wSvwWRPnUfmFnO
C1N18go8LOXNHsqQ8igxLfOPcRELdM8fjwpzwOIRdmcBUsD7weesL9DvejjnqQ4Z7HLw5Q+AEXRU
Y+5l5NZONMsHTGkx5Y/4QopP3g+k4HOVDP5PMSG5u0Ck+Tes46ZbOmVuWw5nWsocInHyKV07UGqs
kaM3w51rMog5XJBqXDwq1MXkdSnwHexmWMzjVWPInh84OshwX3/p+/IHbIhWRl2iv3QIubgBpT4U
OI6SaWprUkUsE41ueq+NRhVlvXSVG9eQX7I/GQxeBOsipPjgFp/UqrD5V+yZ+MpzOEInpZn3/ViU
R+V8lXqu96MsKt/k/IgQAS36iSMKNlKbggAzEpyt0prN2MTMouMpWnOjTjCfTWksB72J6HleKMyG
sRj5KN5LcsYz/d7BS8kpv/FO/UtgPTlZl25iKcmJhy0yGlAFsK9e3Nrx+lob/fMqIIoKqCBfXJIK
E8HrJ1t+Dy4Xz/1wMu5dq11c++/rn63pG8FAXIiZ9Zp0epebPo8fJmGDjly/5RdJ1dcaJnoKZ5Iz
XWHqW4Xr1WnUuXyvBw6vXzhiOrVTDMEEqgPV2+ixeosjZ3xVflVfjckki/aEA55qcqOPd7tBSWuE
gp4sldbO980TLMVRiGDUsXlHZv2g9HBidqpPKfryk9J0PYh+mDj6zqmHMl9/hVrMqMOcoSLpHrIs
YJ1NZjRHs+xEOT/hJhehof3MD0M5qS5QYF7XHxzQfJWx4sjoYMIv3BQL42bnk980ZNzi0zbao4eu
tEQz3IxFh+czbS0KnW9kI6vh2hA9A6NRVR+0wdWjJks2+LeWM2KvHnqxKyl32KyA2p9u+5eh/jSL
mrjoNLLP9L1ahbiXCUtoaUdVnUoeTzngcFsnavTBBhZ0w+fcRGbU0k8pZZpU7PwSTDipS9KFCi1F
pZP3EdSaITVSjOpUMpcpLUCj30Oyw2ybneN4tkQ7hGtSHri0GSmNuQgmC+OqUMoNNj37GwAqgLSK
cTfprGR8w+M5qvbsbmHBOBGXSTT51s2HU9Bd6hDgquH8F/MzoKLR+1N/3vKAg4UK5bOZW3LfqymT
mHkx8M8XR+iO4/70qnenVKSH3TLa2X7Q7qTzVVyoqQceebKHJGHK3NfgKl7Qqed73daSECDTFY0F
o1BURKgwHSrFK680bS2VXebBI7cX/XiCYguBx8UueH+EUUE4o2EXNCjzuoYReHjdQUFqssSULSBn
swGLLl3i1sgkFbnYhvQkfJmKPdhj9rGbyfns+iwa0+uv5yOH0iulaU7xKUaiO9ceFWhIfEm7vIlK
xKNRoztXLKPUjybYM9cDJNzQPdNgFg+CcLMxnULDfWwXpfvSe9J00lyBceaH3vBeSuyKB+EwUeRX
axplRPse1x9amg16v5TzXK2CmDZkf1b1bsVve/DJ7Y8A14oqmbcDBERj8oiHe8Tg7fEEnsqGdTJT
OCKgsNEsuvgm0ZVGFMmRJP7KlDHJnVEMcENdMjAXV41sOuh4qLIg4vRk0mF7Vnp8ZE1bvmlclHPQ
H2/cdv4eYsOFieENawtnO04RUSBPYhvGKK70KNTPYfP9CYVsuYX54qOxkZ6WtVOWGyvruDCi2zFM
muGiC0NpA205KDLqnDdX9STn/humomkgIO6Vy2/sS61S2AAgWw1HdHUckuJmMvSDf3+9Uz4rKYFr
Kwb9kMOEUbuBNMrhTB3MI0RMmCwQ6G6uHJATkuOIOZZ0hJ4VrsA2rqkC4RtFYYu6VZHz0GBoQiIm
Smkz1sjlykaSdZmgrIn4ul9ByXBa9XWXoEneGmrrBhhIy4Ri/7HqtpE7tDGbyXrNhg/MWFrNKvWN
yCwqDJTwS/wV1pAvaA79cjNNXLi+IGff3ixDcilGSeRZwlRacc2h9a7z8m+ZdIX2B8ZK3MtcdHhP
jnyXUW5uXLjyByntBq0vVeKhFOFiVer8vOJeyLWLM6xQOELRDUq07Jin3MGaRBkF3qifYETN2pSu
6h1dIgAy2rPQqtZukf5ozXZFD0TWCkYvtr1Qtli73daNlvW3KUnPQ5b5uwyLShc3ArnPgSDwVr96
00eXkO0jYAH4fV3Hgq3ClC5O5hvh1ZBHLy+x5HInGM8SOgH/a8kH1KO1hPW6ruBw2i61Ul9ywPrT
jjPtfOkslV9c8Vns8ilvFTHS53cUtE00Tq+D74Cp5NAD+440GAW600FBa7BkJbPUwxVWiRr+H+X/
2V8v5NLdLQYeSnA1hGharmktn/ihaxp6zM/KsJovFHJPiObMz8EOLuiC2sKAq4+X9iSCbCoTHMu2
Z3eAhQjKsTEoFmBu0JdHtwKi+1AYkDWRvmM4km4R5N0hmmLqPUJyAmG6C89QCx9SVWRMkwOuCzgP
KPEQ4oMAfWTEVZmh0/kpOItGUC3PSrbdVdEYKRQdmGGNwCBbKa1no9eaJ3oCSR8JlaQbA+0hNxoJ
c7frpQlsutF+A6P7j1NM5biDrCozzPBs51fSLuXm9eqCzjTCvbmiT2+dNtpuu+sRPR5M6Kz5hfLM
v8L+5eWsi9keP5gxWfhjpsj9MnTp4ckEIg407a7n2BEj3ihrplXlBsdW+4wRfOV/BMBb+y+dGF1W
kgpywnfgT3/u0QnJA+FkMoVvBro6t71NuB1zZCisB+0jDEKPe4t3ywdQN0hTO8wPCSb0XABpBWnc
4BGVHzqUXSwSY1fUDN28FTGHL/nAipdJDfIuEZm78qFOVQvMB47l8xqH+a6m322XERG619esd6GZ
4kFbcxkaW3hSaeAsdRpDlfkm29C23Vp5FzyipFoQBbFktOiWMljEtpisQL4x1K0zrDlg8XeWS3Q8
sX/tBjJJe7F4paoh8KKXLoz/053JUREjL92SsM8PVmcACbycOJp7FxAa5TlPQfkz/AEjfYXPeJ5V
d7fB44MC+HkVbtSnbcHIu1UPw77I3YNY5+F4SlM7LoL1cmOYflEpUBdVXZRRagRd4q9+uJ2PG5ZO
YkWgfuo4OoEjjHyDTOQUo3fPH49rudOdCuFvw310VUm7IZsRocd0MV/5M2ix5gWxBv8fe5P3EAcJ
/jWgF6JdmZ2y37Dvuu4qQbPF8cARlZAyfFkeBdlh/+R0juTgNkifhUEN39K3b3dL4Il5yNzjyfVE
S2MCO7SSSWFEuTu8l/0XDwfjd/oB+rojYdn+iuZTBMs8pMYEpP94Nn3ckJL/cql1wa2559jzpsOn
Zq9rWJe96P0B7SvcD71WFTYMsrK4Mp7h4R0TSbqaw6jStX8zcMXY88EgMGxPyY9mV1EWTD3/HXGC
zIvWPWmobBKcoWG4QNr0q09WDrhrZRLamZkinV764rKymOUIObQ2uUhwTgc5TSwYjeJhXcSOPP6k
nf10N7JFsXdolsoXbDS3gAmShHBWe/TTzGtjOwiee6nnQgT4KYMX6+brLBvvnLovmbBvxNsaCIc/
ljwnqRInyjqZTzIlBdWJIPqxoBAWaORup3sI/hsEH/srpIvwQ7OlkPlu6yk9uf7aH2cPU3tngdru
QEcxdCEQwSCgEo7UA9bpFm6lepApBDc7H79gUWNm9WRz2FyCXxzFTjZAmhb5z0CDfH545r25kx3w
4s905YctQZrwiE+58v6ArNUavyNoa9HBI0T5aevLNnI93eFJpLH7EW4Xe4yEyzyTCEADoiAon4m2
nXuqBjzTnjiLueB8MU1fH7S5+oZVtE3Q26mz4D3ywYy97ew5OFt58/S4zr7Ep8S9N7rzAF5e+kUW
QBRRC7HTilQSo8HL1MCO8SdJUWfkc+m5yEDh2rAKpD9IC5yMbfqQz7uUDYAHqfKoQc30eE6J74Qy
YPrc1MmIYx6qmuXYPmvS+LZbQkt3iOfD0X9a2sVRREQFDhysA6sCR8yFT7D/t4hZcfAEGWpWiqk+
Ln6aM64DfT1H6YUdr15Zs9OHCZqbjlRB8uyVTAN6N0u1j/kBKPlt9izIC99luSK85v+5l0F7+5+F
BLfsQwecjDqkKtPxNCp7cyLciX86tID4EkS+OBs49lnU67C1ChFDPIZfl9SnRzYfbA2107780Emz
9PFl5u82MkPVTu8p1QBLo0dMC70JCHyfrlQjMOCi/2arnEVcLdhfibN6kC0wrdb7NfI2OdWAF6Uh
jZdj0l0QmOwKG/iWPtvkrMSeDyybJNuBdf5dXN6RRzE2cdjzjCAAdSx4x5iWs173iWNmtAp16goo
G6d/3meurAA867C/8c3j9D+vLWanlchOk4OQ8AVKu3ggOHSChIgwA0SHCEKKBvHho4Zfn3Mv37DI
WcYs6lUtZZYPzzebVs6d2Sab3+IhdData39C8hkI3cv1kWNJclcQCn5jerxpfWGxfiC97lCTm7H0
ePwW47ZjwsSTncEUMw8xFlHCQ6nu74GnNLALoovMtUS7aeaakdQTjaI0n+yChj3lotD7b4k+Gksw
L+PStc/2HUOAX2wqNREkXzwUPJd7V1fKpBeL+X/gCauBeA6jgDk57Kh9T7BllQpP54Uc3jeko9m+
HGqaYpPY5xbs43v3s8mihob7RCQZPm3dLc67BWWVkzSTDlOSSwSS8g26nzdPWsRb4BF/kke6x8WC
b7OGlsMdDU/apySdJphA2zkDdK1A3qZWQCmY9C2xFRA7yXKpaqKtdCHPXhA42NnH9AfD+2pr30dp
iFPOVI6i6nrKCbAPe873XkZAmdd0z6zdGejex8ptNCYwE492+/K0Sr5EMkqX73hB/+8s2Gj1sfa9
1NGLLLVjKo2Ax6fURBcP3Ctrp6Md4GgL1Sr1WPMc7BJyGSH5KW7yDIbTZqZWsfLLgCQ3OBD8ZW12
yx2/PRiCGBX63UJ18Qq/VH/NE/+036qiBV9jEy23n7CXXX07oyv9/jjxTLpWjo7utUkNYD7Y2uTU
e2ZW2InGpT3LycrQxTkY/eIXOOInotjklT56eNbsgbByg/Jnb9U+KlDlDG8ruKwzY32Q2e+l7evu
etEBbg5h9RjMsRdEckuv0hZ6en2EKKXHcDuN98vzL4fKAssXCZP0oSKKbpdsodPfiTdm4H5xxTSl
esttvkXr5Z4/bZnz3XUSrX3gtOUEcxOzV7VlhH0w00ECP3XcYtkyK85d9dgLatayJAZsvYpu7d1j
yQtx/yRhoI1EJukETGG7kucChqzOQmiQ2Bgloky8SQ+y3Ye0yO0sRTVjd306snmBcvnU8PxVPGux
mixEs0JKxP6IOUeZLKwlRWH9zI5a+iHVa1C6MqOHyZ24xDG1ePfMX0g+0CL1z6YyaTnJrFZpdY6C
VXiJwOLvhyRI/Ar9acmn145IARWUpJHdtrXeRPpwQkCdRVPRNmLAvUFenKujT30RXEMZ+hxAIgoo
rg3HcR8L0nGBfzDujheafpkdsebQ8XUMYuDQLlX7jck0sKtEl8c84f2ktT1hSzIM+2UmLJ+RZSGF
ftSw1TUi8T+pZlqhcDpesroJZQTKL2IAQqWpLT9rCRpa7v9HtMYuW3N/KD/jDLsXOkHCoyMoCPBa
m7CwrA3m/kXgvPWyfJbtq6ylINFPRn5vd1tKka4Ol0+92ib31rRMGYnY5l5yEmsKOkD7KyeN/Ill
nFHIOTt6bxNJZfWUqlLdJ/izvD4ujlIj+3qrIvEyp/TPZdXrFxz5WwP00oub/B0greBao9EtT6Kg
BZWylqtyz99H/Edcx71hTpRC5sf7Txof+VEHU2vM0QkuzTOCiBDkgVOV0BC+XqzUx2g40/tIAS34
v/D/hy1h8IbNIAPZdtZ1bChW7S6S5sFUQvwqvqNYdnD0DgW0L/lidYcqQvpsCCMjnC8fKcq/JIrm
MWZnqzAsL2ck3CyZxgOpm+i2+zy5rj7FpFcgpmsd/sYjdAxvK9hvtzE1vPC9t3OXhwQ+hzuNmiUL
bSg7krUoTvJQNt576NuznI1iy01/pYDE3zuAUh4tzGb1Kbmm0rDfCdpN+4i2CHFbwgmNCUROSLw5
IxqqAisEi9WzLEYAVGD/dgs4fGa/Bjat87AMVYW0glwvNeIqw9y0vkWdMv0q1CNd8BSXdhFbmBtX
UtCnCq5ap+Gnz0u2UidDkvFjlgJi6pVWmvlzkF7zXAF3d5XM5eqiB98CfO/+Cp77x5x+JFerVP44
xokqhBL+KkUMk5eFW+y43bfpF4DB/NaIWb/EIB2tqqZcMeKLqMLiqJO1xyFxiA3yEaXus9py9ebH
0dHYA0g66ULDpKQ5iZze0OnEM6DWFc7Mbarb3IjV9IYS1HmrqpkquTzk+HjkfRSk0mGUQk1Dj1XV
PklXpcKciscXtSuxkpnU4uOuDX9WfZj+ZTEUKutcUfhoeUSDmqLwgDnSkAP4dyj2moohluM8dxeD
GtBNyqSwUSJ4Z4esm0qYfrMJKsE67wieIp0q7JjGeVDZWu1LgXWJxPGD4C7EM2Ff6Yce1jI1AzrJ
qGKmrqygFHQXs5VwhG9INzToRuzOh6LThxEPu8/aH61YxybaE24Uw+NiazlgDdFppHRTjNnvHJ5R
EaabNsKb21jWAIs6xC2+3xs5IJLh/YaqX/6plzZ1NVKe3mPJUIk8zb6m9FzbGb98hmkVKQZ41k9i
PwUZ4L36z7WUHZvWrn1+kjvTbw9Fn8e9Jc1n7dEcaKZrkeCqPC80wYu4QbMi6ZWWpsUrDJpX3DW7
3nAiEBMHBvySlalPZcY8XlAgkBcJelbFTKSYsdEm53d0k6cmlB5cbNZi2D9BSA34kUyKmqIS10xj
XnwyHd7tg6qj8Q6JzkM3+Ybp2hXcou9hHe0NWA5rcWCP0PRYtVTeDRlpoTXv8jCzVtoD9yDFt8da
/UbXf/kHZjeOAL0bdEn0U0iakeqj//J7lMHi6rOsnAVaFRgXQsFrOHI9zvEhE+rR9qCBzPoO4sJt
NoyEHYnox4f2ZnqoERpNjR89wrCNngGCNBNh6rwwfyxv7VdNIIaQaol2XIg37FA4qe+NEvya8yBY
A+TMzqhuG0VSGkDfB3RNemyi1ZI+/mF2czpQbG6eaGpqp/YV+QnuyPusNrXUlGjArZVsMDHl6aa0
4MDvMKV5NoO6rKEM2pnYxKSppi4hWPiz03MfBrTaVJvwSzn+oy8u5q2xySsuVDer7+c6+r///HOe
b61XrIoirFOfIyS1ODAHw62bMUX8z31l3W2XBPLH2K5b4NqAb7pWXO4T3P/2y7OxGwBMAQEztcsn
ZAa31gYIA1IDaXcWv5K1QXKoIbuGF5PF2in8KxMZVHc6yC0XJik3c5oDoynexiM9JwYu5f6NP5y4
SwRextM7m6oYMwZ43jXTNiTbAqv0mWBILUJ0ext36aaeadhrOtaRGUZzx+Xb2UzX5c/LYNuNbNee
fsf3ro0L1R/1+NWgU3McVP+inX25q82s8XUdJ9zThBM3sEA7KfDDqimfajGk9GaY5Yn0XGx14fdK
tfBa2xHmMoMKKBvE4/yjOabItc8eXogdugsaiMAgGffTGhaFWYIBrZ45f6OaZlMR9pFOaN8Pz8a3
KGHvNe+Sul1OJxRIClh0JS5Pj8T513oLAth7m2XPmsT16Yzbm/IG13xivnJ/1IeMDqW+zLPDfkto
E6YH9vovfC9RlDXP5LMy0WKKfkTND1tonK5LKBLPoQt+LeCL4QZqXAprhFljuU4i3/uXCwoHB4J/
ceEVOdTDr2CYqhUMxYZC5Ag6/8I/44qSwyEzpkwN71TygyBk5FZIoVWCkwsBDVES3Yy4skqoj29j
EfAYIlkDCIuO5OCykPAIpAmS7ZXnqQu9zQp34XJtxbgBAcyA78Wgg5WWoZ0EMoSZHXHAVLysJLKP
if7NWHsz32BRoD8xdJ1WaSS1ImAtqYPOzmCR4BwasiijeWyhMfrbIkljCrAlvvzogdmD5VZI4idl
nIoafN3M+fyCKtTKx7njjhwNRnE7QfvxpQS3WdN8yadRmD30TEIvMk8AHuAlNqXXFTn4uBfBN9oR
WRP50daBN8IJkENn9hyB7xo8rFUhcgsYFAFV2HWxUGpGxTtRt83R0tBmGAf1a1w6F1VtirCA6wEg
sg1TFDLdnz0Bx3MPOVqWKZGFrGUE3Stg9So8NhUGD+Jb8pgEvNTaRFs1ujnwINchE/T+z6bYzgX7
+t8RhhlCN3JKfy3L1CUuUc/i9AfTohXzazmICn0ycbtAYGhuHeLp7klPPAyVTtNwsHMprxXnka82
ywCXEw4qdNJeCYv3Sk1BzyMoLAe34HC46QutXyfOsxgt1VQOTU4rCyt8K8ZxizsaiPLY+b16JFSg
VgROABIPqYXdDCuMsybjQ4ejOZNXf5a1dfUWDELQVGkYR7DJsfuky/+58yIACfjTWT5iAnBrd6EV
U22RFarn0Gq9fdTwPI+iefdrrKAI3B2kwKPvcFT/D4oimUYblVLBnXR3KuZQEM+o9ipPdXvVTMOK
Gg91/R/H8pvDbhtp2oQjlzGKGJYQUbKIszA649a1IAmHqy+NpVt3/uA8guZCnI53cEM3PbH/orEZ
FD1HMKoJNyi8sgcSxKYyS/RLn7C53f6sUnqVJIXS9fsPlljKee4BeJkvVsgI7R6F90lmImvShj0g
7sGz9OnLOOGNlcN2g6d8Av8k/yHqBcHQGs3dKINn+F9rNYeEI/6PPS6I0P/IDtm2Pfs4RCRcQxlJ
jIwyUQPsyyqVGDyDKZRc04Jw1ICOrp27JV/xl54qySd3pQXl0/zUlrkW56l3hsoJQWEazD7d8bVQ
vzYJRSprvboQ/6t3U5GctT7hkxGzmUOPngVePhFyl6gspXEb9jLSMOgYwwFAx+C8TeAPYduyfdvC
SdnwA7BSQBQT9JoyQCVNERoKwGOSeehkEZefaTVNGl70K2zyMSFvFHnqEL5txAxu/hge5s7F244l
NlHl5FeXBJtzGHVA5D3Hu9dlQ0FDh5bTRyaJ9WZOjqUA0ecM2Rk0CFUob4WltBgpTtZfH7F8zZJU
EDYs8joP4eD7yRUnldgQ+bkb/zcDxNECAYoYOV5Z+98fNxlQHdNA57I6AsD8gJ2oOLWAUkIP1TMG
UzkmTkyD/vkOoUDeEgm375e7l/S/eo8I0jtPcs0TzXQmvlOcXH8AwJk+yYO7Yk0vtcjqYsMzKm9G
iHxX/twI3qLvuJT8iwoLno8IaOPUCFou4zlAjwIvJVG1DePvDCO5G/5W3HJjjX6X524d2CTvy5pA
c7zqQ3lrsfjxPyvvBfeKAtv33QfvquC74nDuL1ttEFzvgFivQtau36dSw7+vUtiNMiVvos1JF6Il
H0/EAR/GLw5p3KCYyBuaxJVwr6qQgPnpIK2omSf3XiYldKq1SXhMio1lw7wfA1oekjgWWrmFhyLw
INjm8/hTcy9mWZfr5Cj+6vN9G5EpqdBQWkcXJcKnZvdwem5DMFDQc7LHT2K+RUDg+Q3Z3BVFFqu2
m9rTFDGyBz+OctGv0gD9m8XM/8ZSbaL9vMON52mvNB7qeO+9GTlLvvP7Lt+ENyHil3j5RD2BfIzZ
+tFcSQ2GAQUM+mgD7UrQ3UdS9M/taFmaEuGSCaMOIcewaRtn5CbGEaw2gVlrcP4pOTYQSJbtlQ9r
IAV8q1dMrLcMcTxL8yrCMegHCsW4LQsz4FbAF0TOt5HPmwNaiksoaeFV1bobV0RfHxsXpglV3/LF
GX3QzFsV95vWFegiEyCMZ+abOs9tQp6wh99RzjeW4kE1UkbcqLlgLZqbw8sxEEm3P+gfnTx0611C
xBgjot1CNCwVQTJer3mLtL8mf0XYLVsMmxrb2beI6XYnMZakHyfXpl8tXYqO1AcKpru3ql3F3P2x
3SsvH8+QSnl9lH7aBzLs7MQ2MJvga2hw5UO4LHtDZL04EUPQk6+AV+3jlFMrKNZEaaCYbIAveSyV
3blXk0M71q6f7Wco2Z4YHNoqOFO9oYruepdYWeJNU4GeBLZ9Hh/bpaIEZMOrkVCm7aRXeCtyFG7c
UlisdiekYML0n8ShyXGOkJQkIx6ORBNBEo2AVeYSbzV3cyV7utUmwVEoJObVq2ONGkfYCtb+QUbg
Pc9ApwXexBNAsZ1jF4GnKjJ/45TLQMK7tz9Ql/6roROUg14GfZ5tDJ/oUqOYJPW3hpk6wcwUCFzd
zYrA1rxIqElinkorsyd/NBBsXoP5v0eaN9Jdr0mWB10smUoRJoLVhNawA03GCDKCdQIx+od86n+z
egxyUkDGFe62yjFSFB/RqidQY2yvm1y02mExf4fOu89IZY5dUlr5B7HVgKnNV1Au6BwxfCpdU33h
gS19f+z1WR/IizcY+FKz3E/5Xu2xjfvL4oWoVZlpTrG4a52IxVywwZMRGhr31oPPo461uMZfhDE9
RtSyxqNWUdz9Xhqogbh6uAc8v9rwcs8HuyJPq9QL5zf5tsUgA0zBVJBpzl1HkD71+C1zpFeHIt5q
DjNH4ghI/v+uIrfj4GJVZv4mH6+ALpE8ZIkejhiEHa90PHH89lHwOD4WZqNAuHf1yLiZRbeSODrt
MZxgleBPJ8IvsnIKsDqvlyRsHSy8vFQUmFtPqc5KFnLFFdVvmS/fM/kn1c0gghnX/xQvbzIaAhRW
tMKv3clTjX2ydSANmFy3Xr0aNra+M9PohSPUY+srsM7eO1cHr93Wmc8tdfqQF01d3g9kq8paBQGh
aclo9V5uSqDFODYzMZ6nl1RxCiVXVWCU8jhmXm71i+3tzup0yeSsGmKqbHaoxadxb7eBQzOOQEvk
2GN5KRkPzWPl7h0HJTfUxp+yKeo/InP40eerJ67kY7KJIfTNAMWDGyqgIBYZIPVWxuUVUVfGpJN6
1xsk10ggoSIl9bWiHCIcZKCeqkzDPYvJdOAUiGaK2hbEBhHVaiOC3+QlzND2VcTiAGNSdK1wxv3K
zI3v0eWVQmcVVjqErjYoOHK5Pme1QVucn+nuhimlFIS90mBah/3oL/7NIcBiHYZg95Ldfr5pPAaK
Bi1QKWuIdJWm7/oy2HieevFYaq+Z+WSa/U3hV1kw7jNrNi99Pf+kSRy9WLlLsmxxjGRt6qoa1pqv
8bn59CCpB3k1Da81NvZ0SLsFOXDuxz1uD7ShemNaeMt4QJOab26ihgkEmg9NJgk0zpQ5m6LuBuKi
8eS08q4OMSdOZVAWn//nGWoC+ppRAWT7G0QOePj7bt4pvwGWmxbgzPZ5mcB3KrDkjYb9UlTyXxoL
rRDaH4dmCQxiP1gy1aNMyD7DRtNLtPuZSbbwwvaIRQ4dO7+z+vv3l6p88gLHc0FusJ0jsVeUvWa5
+NskjUGEa+11/lEyISFeFrG9Mct7VthspaI9ri+f0qFYS4Bm1CneS2VOCOOjb0nJZWoOiXhT2Wl9
1FrL+fhmkjaj/pRi7Hgs4WcZ3ft9H19unXOnM1Hhcm/zO9YBYsC81O9vUgAtQ1fmoaWfhRcUnmvj
XgAv/FQ9uz0CH1w7B7QMZCCZMqE4K4sOMvaxiLpeFaim+C/p/pcggsypfvzqaKR2cIdNIVBTdsgF
RHHNwTfXQLRUVY0Hc+sBnferp3dNXdELHhGHUGlUp+p1bP17IlZIBr+wY0yJJ+4XM3Hgq3fIsqcv
RyUELo4UdgnS5XoIlRMqZ62lbOOcoRhFDDy0m5UhnClnEqfHdSKZ7XhQb++33HsBo3yK1GpwUo2z
3yjFRGJO7gTPy08/2+Vl0k8F+SbeOycixci5GMBl5gzDQ+/qDlnhbQbX5BL0RgM8zqOT92wsj0kD
nzJYtqnbTWJPnyj05+F5MXINELHJaglqvGWL7lAMS7x54s89dH6JEdrDLFaxB9M9IfRAcLZGtPRZ
r0caF6deL/fJeFy05Gmp6h0wuNhx2Cej9frmlm1qFOlyls88rYF4jgzCyu8gpGbFKhDjtigiaOtz
rO0vfZutf4h5Cu0l7kF8T1oHRWF3RI2hs8GyGb5wMNo/Y7JHeOWC+3iRVGiuOc/7StUuIB3SnZa9
AxJS0r1VwIsiYGVBqbJ9KlUOyfXdlqHsnpyYIkLsReBAxfZ0n1c1McEB0OV1aDr32ZHal9sEIUig
j0jPZ3KlO9BQvH7dPUtRhGLCu9z+bBdV1VUXqs8OxkPq51Qb4jCuHdUlNjSWjD/gsjHav6UWdr7m
7hU6FCkpqAtrlObSOJJo/VN69g27+Lt9658pn3vwPBb69R1NYuRvlGZ0xhmQicbA2S59ncIOQ4Jb
U92uMALtEZTQeNLzdAuYiX8oUJa80hOJ79vm4/JPGPQs81fgA1+xAkmGXfgwMVWSVU9be03kfllT
q+e8V7gfkycEPhpMH1wT9mk3wUwRGKAPL/XRdawnW1OTY4/8OSIbKYgSDv1MklmiV3sXFryNAM3I
p2QMoqNiT494v5IH+cB2RTrSGUl0gNQhHetY6raRBpOY19lTXsF55pXyijCOBJtSp668dcXPBkTy
oBSP2HpWWNdeypKHvyItMp9FJuwXqOQIoKSavt7RH82ygYUinRHf/SHrSWfY/qxP0P4D8VwQyifc
D7V0xc4T5jdXFROWmct3pV4q3gOcaxXn9VxaxqaKbjhlijP8pRvLv8caBiyIx2IvRDX2SnupA0Mq
I0JgwW5AybsRz5zKqm0MCKb5wyP6bfczOQKc53sTt81c6wMkye6dnEEH7ReMF6Asqm78dSzZdE9b
HV41lYCZG8XB68Qy+IQh7coKWcm2tYetf1wWzTk0xUrCob2cMXX8oEZYnA9wmcW8QpF5AwFOoK4S
6zQcr094e3v2Jh2gzhMWOC3D05k/8RZz7cHtmP0yi+4lLtrOLgpr9STMiPYEnLoG0vfa1JTxbIFA
eKC/THalIAGnxjoANNIp6QuiC+DbpV9dbL4f5W+OUV6tt8KEd/MQ+dpZR44o0dYjxiJjG6Pf9uHi
f/+7VV7UBt0xJhEhm2F7L+3fWWLkOZCDEhTD1eLRm15nyj785aDVRxC3wQhoLqWLvTxNEXKHxhte
weBReuOazzi8LTgiFHzDJtB9wFN1p+25JUAl/82wwrxhf9L+iK6NSDqleZtFfbc1DR3aTHhccn3W
HBwQmgEfdj9fX9QB1xLmPFZb8ciXENsh1Op7hUuOovmotKDJ2meF9XLc4/0U1jJUdNHNvBIblTIU
LIR7ddWHTCxfLnqT/uMQ/oz+pzNGV6z0rq689Nl0pH6tU9wTPPEeYuA2o5DVKiwXx8leUSb8Xp3R
jP0XN4WS40KbUNadrTTyyf2coaqKxXe990GQn/VkdfNn4yuzNsXYzWXOMj4ioSwL77A3+boeeXfo
1Ru2QBNAALp0TpwHbT21QBzD+E5otXqBhuu97qcBRhGQRXaaAQ5pRj8X49ET5GKUqyM0pW9iflP9
nh1WhAYgIp8IY+DWor2Yh+i+B9RGJwBwSOEJ2Y2AsAtwp7Ss7IAv833dQcnxsMHdtWc/KKlo8kb9
SWCIlf656/Z1OofiAlVG9VcDWE9rNp4FbG4goqSzGT9RK/o4uvjdqti3FYnj+hlUH/gQHbSPpKYT
OXV8gae5IgIFRvoEpscgfcWb3ghpP4TLyWMbj0OCG/4a5KzioBjOTivEmikYiU4moFS1xQnAISJf
KGwbvNR3tjn+tT7H0C0x/dD7roLlf7KuVBiKI2eslFK5uoF6gIV5OlrRADxV52L0Lt+j+SrfYfTC
nA2OPPysTcBr/h3Xq/rAB1P08f5GfSrU+UFcY0bpHvt5CFE7UwpqBZ7TxWw6qUC04HsB0+tLE6Al
v1b3bpZ8lnxvp18Y6V43dLRD+SGNzC7RCEVj9CMYQQoDtFROI7jyggGVYtTSHMxp0pkTE8SQZrJQ
ZMXZy4NXVd+Jzowgb6t61Ukd542EzTIUvrnMRyf5gGye+wcc8GX7jYQJWJqyEdo00/+oe/LNGo3n
qdSlP/22Gi+uY6iNJqJrXR2L1aOjhuSMGQdkzYMWzrNbb+fpjgxkQE9Q+yx92gNUoYxPGyZUd/La
OVGGyRy62f/61E45XtTrS24XeCXA5KsEMWiYUiHej0H8Q9wP+yleAHNOCi9SWp0jIbLmzDI3c6+p
lRoIPFQhjxiiBkH9mwp1eb7DhO1AfoxcaFK4AZSjWaPAhavzMH3wzO9bXfivuQTIJCKwpi7Ne3js
4IdjfnEevLzNTBt1qzNauEuun3j+7cBigDjju3xwZhsYX/pzhDwbT0KrJ666Io2IkoGWLkLBKzcV
ILn9gH/zsy20ZHdQzt/6k+Di4A4yMOxT3ujAXMQLKOz3cCPSxAUYSbrnwcB27Hc6jhfrxPoGKkQr
yecfY/uZv60p6tH4tUfwhjzuSuQbNxjzHFo9HMebbyzCj0aOc/NFrcx6OmiviwXfFII+Ci+2TA9q
lNxtoKAJG3Eo0Vhrf9gV6uV8zehh1ACEUGNUXKldf5CiTOS2gOgNTHw4ht8TAv+354rQ2DCj5dGY
LrB7zl39cN6q1JVDsVobR7Dnq1jx00/Rn8lGjsPesD+mSXfgW7BrhPxHcNBCK0ujbL4gIMIe3iFk
1bv1IQ2UiAs7hKouOm3YIS0B5/paLX94l6uYbFTbzDGqojanFFHNbSt6iJlVEucXZwSGjvT2q2pp
NWlgRwTHHrP6EMBpyKgeAdE7sUSQEcmXxnvyVg3LtRpIURan04zrJaBtZiUaazgTo08I5xnVgL8Y
/SPbc1cVt5Y4AgcqMYBdxtFPWbU4MPf8MSLTzT6OM4k9pYZOZrIlQ8ITcIEYD13/YN7ttO9ho5po
bdj8kiQoIWSHwZqZr+6/JVcxZ2JU+KgitX4Yf1skaUvr4my4E1GcRw6Gw+vFVO/k58SRcjtrAlUQ
5JnCnjwoBfoknA1BxNR5DmwhHv9zmJ/KTe4+1oSwnZP2FHJU9tUAal9LNcnYF+lCB+c1XREOa+WF
FwP4i6sptGs7XHaMtulbahLF+peENVunJZ1jrB8g4Yi15Ae0dR1bc4l8ldKy1l68tAh4eX93j5Xo
Xfqc0zIWiB2lnLAoNWbYQouQrLLqfjhOTJ1T5EkeCGX4h9e3ay+QD9Zurbp1EmW+MW50M0tTUZYn
jGZcgXzf3ECCMv7QFtqLKmUd0bP0RY1c4oFTRcohogf5xhL17c7iiZnrkMAymNIL3B/3gYiT3Rv2
xddKlE+oKf+cGYs5rLXhAWoI3QZAnMr9A58wbdZQbmi2mjN8sgtBinRhe9zgbskn/7TI/hxBEjbZ
Ux4YmP2s1R9YzPp64ryuPyAJMfsSG1rwCc1SqclbqnvxSs6zFa30WNa8nurfj4fTkr2jkGLb8QGE
7fnRz2AjT1Og9XL9oPfoWWdbUs4VVZ6YJZIAIhpp8zRScxKNqkGJ56GmQKYYnxxCXAX2A63cDNzw
Kao5DSiv7rdIr3YhGqQisGg7MuRg52M+qvi7JC8L1LKMRky4eNY07TaAtv1VoM0XaTeabew/sU0m
Im6dUVAXcwJtSfPbWvxvLqIO/ttLuXLevZI/CnY5EnZEBjhWa4LPc4QaiTKZjVSFPZADHXhH9Rmx
33U5F7pf0ik8W4bl36vx5vvUReiQwTIfcdZEGTehgMS5mQwEGCYm857dWco+wfGFTrWMt/izrO/V
BVuNnDMgZ9PJPlP/9ehVrH8jvMvoDyAOUjgqJ6ql3tiCJOm+uJERl+bI8wv13k6hRgGHY9RX0n0+
K7kIdzwdF8qAzB4LN3bmfILxI8NhQxucGZzKROL0PIqSsnS0QgAhGb7Rv2lM08SFdeRMOnVaqDaf
itIWFU70DtgvGEYIUFFZew22t3tvnnomvkSjJlAe8T9kZS/vSvBeyq9j+819SqyL6vt8BzsbaKZ9
g3AdpD36F9GXKi7MLLeNvRmXKqtdTz/gs9GDzPG68Siy8AfJsvKuDoSWDtCNYRDXWNkqa1zxLwKv
/vImo/6e6MpQeb11s8X0YziDNqupPT+c+Af4xB3WFSJ8T6M7kN+3dj15XZeoVhtaayK7dvcTDSuV
KLAevL2oiRz2pkFVpfcfyZLm2YkagQr4f2htZGOPxJ6Y2UkkgvIaIDpTdRDDDj3u3Q66UJMUYbax
E5cshYRxjaHkAGMDtewS7lcWJSRCe/zeKWcBmf/EaIQwLsBDSX5/0nVXbeehLI/saxhpvon1r8fd
4SjJjrtTs9MNYpd0eAZRf8HVUELvrPJqRYNPtM+bXWm04DH88JtNwFZJT3+2ANo0xT64yEopyo8g
ZeevgniGXaZpd+z845IuH8tUMn5dpDZwIY8OD5PV/kjyan8o7d7/KrBxG6Im2o48YPOfB2MHzwWU
3HXa3gDR2RUqRe4enhMP8MevlJiituW1CTPBLBuwX7grLSjOkp8Zxh1rtWiV83uLW4dANMHWTu7h
kp7mklH2oafFVE3rAvKVpTW5ucJzjJpQH2eF7mtmI6/UJ8wvRGDNpLvW+nm2IZRTckVVMXkJN+vX
tx+IAI+l19HsdVyFx/LerUgqy8zAiSwk5qA4X38VGDXz0QqedOX9ivBs1PAs3Mi9a57bZroGFID6
pYf+ed5uwPr+MpiHKv+i8CPPr1ldQ0R+5X75wNGWMNGMRItFwf7DiZyRCg6W+KcdRkYWVUQJ5kgi
gfuXYpaCYBDPturZoW3sONT+HWwf+ddnVnQgm8DV53FD/1uHZj5whqOPiVfwKT4W9qNU0DBm5CFz
ZJ6NlsVTtA/k6Qji6CYmq3Nwgn+RnHmSXrUAJHI3lIbIQ+ZyEGg82GXsrRXI3QLfv6Rbg6wjbHa4
0FQtKb/RIytH5fxtvo0i4ziO2AfF7uXqrqz214z5RY5REZT9aA7BtUB1qAyRKcbv4qN0pEMC0cwo
ovuspTWWpoOTDoZKQEvDEn6k5QxeQJ1mNpJ1EfGn0BWSIkPAQ15o3TSLS0/1QPQGHTZedqb7ii9s
PFKLkkYsVUytPFmwAZkKr+vCrQpYU3lBsXuh+FyF32Ml/ezueAlCcGCGwlfOvOlG0tNwKwFgZXsB
ZFTbRARUFDoPLdShyO5UnIfBpnQ/NDphj35mYAeKZ/l3xXDz7fR+kCJ+E1NRAEwtBzruQVIwJS9d
ZjE/nEi/W/FXw9lFOv3MKl/MmL9YHoXmXQQHHwddEJ9RH4StEXz05NE7z1eF5hEOJ8RiYsqxF6ym
Ive8hwDLF4aGW3v+PcpNZglBgZ0Wc44G7zfiaoyg2IBAkLi++RGmtCURRjhFM9jXLtrwzc50elxu
faeprJ+WHQRoW3c1V8nitXg8S2qq/aRkEvYJ5l37mkyMi45JxtjYUIO5f304QWRXKVoDtGc04QYA
Q/u9sdBTBIMfvdRPGmzNeAGqUwoJsb1wgN+QNujFPIUvc9tgT9nsN8QYJ3iI5s9MPVk9NvzhqkHF
CdqsKQVZCAPSNQFdLFcpXWQKEz5wOiT60zj45rlOisriW3U1JcjVGX+7qX1klKEbPs0CCtenEdIc
J5WexYpWbDlrQZt/Y9wNGCNM4QZ9n4mVdVZ17fky2uxEwyWORjHaAz7abivATnbk/Glic2InvC3L
hR6ICDH35sMWuRwlUCs9iUEKIridV4wA5T2ZqmkFa45yLuuQBh8hmNDjFn4nKyNqkN3ukCdVXOlT
6gLLxbNocPvP/Nzn6S8dCKGhnUI+VKcMPy9KZy3u7b9DK621O/mTgnr5f4Es7AHtFNVB2gT7teF+
r7o0Pt6CoKpa11R5RV82yHmwz09QI+zP06x/16xn+T4DullWz0TrqszxiV89rAobVIa5sPi2zjKG
+dljNZOvyTcFvG6P/GvcesoTGF77oRR2I4hXz472h3k5S4pvgVaQ0h2JHLx/6tqTnlwIDlf93DG9
9PfXhKyG85Tl+mTFW5sPLWFu81R7sOmplrKcr656bwPKh9Zmn/6jY3So6RYNzcCoTDD93qNVNsLH
e2qKXXAwC5batGeVQmSpZimUz08CKYa92WOJIhgkouQT4HYJajuNg8gBXIi0DNTZ4T7lX+Xqo51y
82Rt005g2jpKcSbycjabvZQ2wkkM1660/Mm3LN3I/5Y2GiJW7I5fM5ZOt4mlrYHv7V2Vma6NB7zp
ehLH8SlaRQI8HOOlm2DqON0RXq8IlxtHPiWyHD2YdM2Egy35rVQy6ftJBl0q
`protect end_protected

